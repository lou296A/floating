

    module v_RAM1_46(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 724;
ram[1] = 1753;
ram[2] = 2782;
ram[3] = 3811;
ram[4] = 16393;
ram[5] = 15360;
ram[6] = 12629;
ram[7] = 8260;
ram[8] = 2624;
ram[9] = 8192;
ram[10] = 36865;
ram[11] = 32770;
ram[12] = 36867;
ram[13] = 0;
ram[14] = 0;
ram[15] = 0;
ram[16] = 0;
ram[17] = 49668;
ram[18] = 52738;
ram[19] = 35840;
ram[20] = 3585;
ram[21] = 3074;
ram[22] = 3288;
ram[32] = 12801;
ram[33] = 35840;
ram[34] = 15362;
ram[35] = 3280;
ram[37] = 1792;
ram[127] = 49775;
ram[255] = 1058;
ram[256] = 32768;
ram[257] = 61440;
ram[258] = 258;
ram[2038] = 198;
ram[2039] = 3274;
ram[2040] = 12801;
ram[2041] = 3790;
ram[2042] = 35840;
ram[2043] = 15362;
ram[2044] = 3278;
ram[2045] = 710;
ram[2046] = 3786;
    end
    endmodule

    
module main (
	clk,
	v_RAM_IN_16_out0,
	v_JMIN_81_out0,
	v_WRITE_EN_102_out0,
	v_RAMADDRESSMUX_123_out0,
	v_JEQZ_155_out0,
	v_BYTE_READY_178_out0,
	v_FLOAT_INST16_190_out0,
	v_RAM_OUT_179_out0,
	v_IR_44_out0,
	v_EXEC2LS_99_out0,
	v_NORMAL_144_out0,
	v_EXEC1LS_154_out0,
	v_JMI_9_out0,
	v_JEQ_109_out0,
	v_JMP_132_out0,
	v_UART_169_out0,
	v_STP_172_out0,
	v_NEXTADD_156_out0);
input clk;
input  [11:0] v_RAMADDRESSMUX_123_out0;
input  [15:0] v_RAM_IN_16_out0;
input v_BYTE_READY_178_out0;
input v_JEQZ_155_out0;
input v_JMIN_81_out0;
input v_WRITE_EN_102_out0;
output  [11:0] v_NEXTADD_156_out0;
output  [15:0] v_IR_44_out0;
output  [15:0] v_RAM_OUT_179_out0;
output v_EXEC1LS_154_out0;
output v_EXEC2LS_99_out0;
output v_FLOAT_INST16_190_out0;
output v_JEQ_109_out0;
output v_JMI_9_out0;
output v_JMP_132_out0;
output v_NORMAL_144_out0;
output v_STP_172_out0;
output v_UART_169_out0;
reg  [11:0] v_REG1_23_out0 = 12'h0;
reg  [15:0] v_IHOLD_REGISTER_51_out0 = 16'h0;
reg v_FF1_148_out0 = 1'b0;
reg v_FF1_176_out0 = 1'b0;
reg v_FF1_2_out0 = 1'b0;
reg v_FF2_8_out0 = 1'b0;
wire  [10:0] v__114_out0;
wire  [11:0] v_A1_128_out0;
wire  [11:0] v_ADDER_IN_174_out0;
wire  [11:0] v_ADRESS_61_out0;
wire  [11:0] v_ADRESS_71_out0;
wire  [11:0] v_A_168_out0;
wire  [11:0] v_C1_66_out0;
wire  [11:0] v_C2_163_out0;
wire  [11:0] v_C_41_out0;
wire  [11:0] v_JUMPADRESS_115_out0;
wire  [11:0] v_JUMPADRESS_126_out0;
wire  [11:0] v_MUX1_165_out0;
wire  [11:0] v_MUX1_64_out0;
wire  [11:0] v_MUX3_149_out0;
wire  [11:0] v_MUX3_98_out0;
wire  [11:0] v_MUX4_79_out0;
wire  [11:0] v_NOUSED_191_out0;
wire  [11:0] v_PC_COUNTER_1_out0;
wire  [11:0] v_PC_COUNTER_NEXT_131_out0;
wire  [11:0] v__135_out0;
wire  [11:0] v__14_out0;
wire  [11:0] v__166_out0;
wire  [15:0] v_IR_134_out0;
wire  [15:0] v_IR_83_out0;
wire  [15:0] v_MUX2_96_out0;
wire  [15:0] v_RAM1_46_out0;
wire  [15:0] v_RAM_OUT_137_out0;
wire  [15:0] v_RAM_OUT_37_out0;
wire  [15:0] v__141_out0;
wire  [1:0] v_D_26_out0;
wire  [1:0] v_Q_30_out0;
wire  [1:0] v__175_out0;
wire  [1:0] v__36_out0;
wire  [1:0] v__86_out0;
wire  [2:0] v__62_out0;
wire  [3:0] v_C1_50_out0;
wire  [3:0] v__135_out1;
wire  [3:0] v__14_out1;
wire  [3:0] v__90_out0;
wire  [4:0] v__120_out0;
wire  [5:0] v__10_out0;
wire  [6:0] v__7_out0;
wire  [7:0] v__140_out0;
wire  [8:0] v__84_out0;
wire  [9:0] v__77_out0;
wire v_A1_128_out1;
wire v_BYTE_READY_129_out0;
wire v_BYTE_READY_158_out0;
wire v_BYTE_READY_85_out0;
wire v_COUT_6_out0;
wire v_EQ10_59_out0;
wire v_EQ11_68_out0;
wire v_EQ1_19_out0;
wire v_EQ1_70_out0;
wire v_EQ2_0_out0;
wire v_EQ3_136_out0;
wire v_EQ3_192_out0;
wire v_EQ4_25_out0;
wire v_EQ5_118_out0;
wire v_EQ6_49_out0;
wire v_EQ7_105_out0;
wire v_EQ8_67_out0;
wire v_EQ9_63_out0;
wire v_EXEC1LS_122_out0;
wire v_EXEC1LS_22_out0;
wire v_EXEC1_130_out0;
wire v_EXEC1_164_out0;
wire v_EXEC2LS_173_out0;
wire v_EXEC2LS_95_out0;
wire v_FLOAT_111_out0;
wire v_FLOAT_138_out0;
wire v_G10_38_out0;
wire v_G10_76_out0;
wire v_G11_189_out0;
wire v_G11_72_out0;
wire v_G11_74_out0;
wire v_G12_113_out0;
wire v_G12_147_out0;
wire v_G12_159_out0;
wire v_G13_133_out0;
wire v_G14_184_out0;
wire v_G14_32_out0;
wire v_G15_43_out0;
wire v_G1_152_out0;
wire v_G1_161_out0;
wire v_G1_177_out0;
wire v_G1_31_out0;
wire v_G2_101_out0;
wire v_G2_121_out0;
wire v_G2_167_out0;
wire v_G2_195_out0;
wire v_G2_78_out0;
wire v_G3_107_out0;
wire v_G3_194_out0;
wire v_G3_48_out0;
wire v_G3_73_out0;
wire v_G3_89_out0;
wire v_G4_117_out0;
wire v_G4_146_out0;
wire v_G4_183_out0;
wire v_G5_157_out0;
wire v_G5_15_out0;
wire v_G5_171_out0;
wire v_G6_65_out0;
wire v_G6_87_out0;
wire v_G7_116_out0;
wire v_G7_35_out0;
wire v_G8_40_out0;
wire v_G8_53_out0;
wire v_G9_34_out0;
wire v_G9_60_out0;
wire v_JEQZ_91_out0;
wire v_JEQ_142_out0;
wire v_JEQ_153_out0;
wire v_JEQ_55_out0;
wire v_JMIN_33_out0;
wire v_JMI_185_out0;
wire v_JMI_47_out0;
wire v_JMI_97_out0;
wire v_JMP_100_out0;
wire v_JMP_143_out0;
wire v_JMP_24_out0;
wire v_JUMP_54_out0;
wire v_NORMAL_13_out0;
wire v_NORMAL_188_out0;
wire v_Q0_27_out0;
wire v_Q1_18_out0;
wire v_STALL_125_out0;
wire v_STALL_145_out0;
wire v_STALL_21_out0;
wire v_STALL_39_out0;
wire v_START_186_out0;
wire v_START_20_out0;
wire v_START_92_out0;
wire v_STP_150_out0;
wire v_STP_151_out0;
wire v_STP_180_out0;
wire v_STP_3_out0;
wire v_SUB_88_out0;
wire v_UART_42_out0;
wire v__103_out0;
wire v__112_out0;
wire v__112_out1;
wire v__119_out0;
wire v__119_out1;
wire v__11_out0;
wire v__12_out0;
wire v__17_out0;
wire v__181_out0;
wire v__187_out0;
wire v__193_out0;
wire v__45_out0;
wire v__4_out0;
wire v__52_out0;
wire v__56_out0;
wire v__93_out0;

always @(posedge clk) v_FF1_2_out0 <= v_BYTE_READY_85_out0;
always @(posedge clk) v_FF2_8_out0 <= v__112_out1;
always @(posedge clk) v_REG1_23_out0 <= v_G12_159_out0 ? v_MUX4_79_out0 : v_REG1_23_out0;
v_RAM1_46 I1 (v_RAM1_46_out0, v_MUX3_98_out0, v_MUX2_96_out0, v_G1_161_out0, clk);
always @(posedge clk) v_IHOLD_REGISTER_51_out0 <= v_NORMAL_13_out0 ? v_RAM_OUT_37_out0 : v_IHOLD_REGISTER_51_out0;
always @(posedge clk) v_FF1_148_out0 <= v_G3_89_out0 ? v_G2_167_out0 : v_FF1_148_out0;
always @(posedge clk) v_FF1_176_out0 <= v__112_out0;
assign v_C2_163_out0 = 12'h7ff;
assign v_C1_66_out0 = 12'h7f6;
assign v_C1_50_out0 = 4'h4;
assign v_C_41_out0 = 12'h1;
assign v_JMIN_33_out0 = v_JMIN_81_out0;
assign v_IR_83_out0 = v_IHOLD_REGISTER_51_out0;
assign v__86_out0 = { v_FF1_176_out0,v_FF2_8_out0 };
assign v_JEQZ_91_out0 = v_JEQZ_155_out0;
assign v_BYTE_READY_129_out0 = v_BYTE_READY_178_out0;
assign v__135_out0 = v_IHOLD_REGISTER_51_out0[11:0];
assign v__135_out1 = v_IHOLD_REGISTER_51_out0[15:4];
assign v_RAM_OUT_137_out0 = v_RAM1_46_out0;
assign v_G2_167_out0 = ! v_FF1_148_out0;
assign v_A_168_out0 = v_C_41_out0;
assign v_FLOAT_INST16_190_out0 = v_FF1_148_out0;
assign v__4_out0 = v_A_168_out0[10:10];
assign v__11_out0 = v_A_168_out0[7:7];
assign v__12_out0 = v_A_168_out0[3:3];
assign v__17_out0 = v_A_168_out0[2:2];
assign v_Q_30_out0 = v__86_out0;
assign v_RAM_OUT_37_out0 = v_RAM_OUT_137_out0;
assign v__45_out0 = v_A_168_out0[11:11];
assign v__52_out0 = v_A_168_out0[5:5];
assign v__56_out0 = v_A_168_out0[8:8];
assign v_EQ10_59_out0 = v__135_out1 == 4'h3;
assign v__93_out0 = v_A_168_out0[1:1];
assign v__103_out0 = v_A_168_out0[4:4];
assign v_IR_134_out0 = v_IR_83_out0;
assign v_BYTE_READY_158_out0 = v_BYTE_READY_129_out0;
assign v_G1_161_out0 = v_WRITE_EN_102_out0 || v_BYTE_READY_129_out0;
assign v_RAM_OUT_179_out0 = v_RAM_OUT_137_out0;
assign v__181_out0 = v_A_168_out0[9:9];
assign v__187_out0 = v_A_168_out0[6:6];
assign v_NOUSED_191_out0 = v__135_out0;
assign v__193_out0 = v_A_168_out0[0:0];
assign v_EQ2_0_out0 = v_Q_30_out0 == 2'h2;
assign v__14_out0 = v_RAM_OUT_37_out0[11:0];
assign v__14_out1 = v_RAM_OUT_37_out0[15:4];
assign v_EQ4_25_out0 = v_Q_30_out0 == 2'h0;
assign v_IR_44_out0 = v_IR_134_out0;
assign v_EQ1_70_out0 = v_Q_30_out0 == 2'h1;
assign v_BYTE_READY_85_out0 = v_BYTE_READY_158_out0;
assign v__119_out0 = v_Q_30_out0[0:0];
assign v__119_out1 = v_Q_30_out0[1:1];
assign v_EQ3_192_out0 = v_Q_30_out0 == 2'h3;
assign v_NORMAL_13_out0 = v_EQ1_70_out0;
assign v_Q1_18_out0 = v__119_out1;
assign v_EQ1_19_out0 = v__14_out1 == 4'h0;
assign v_EXEC1LS_22_out0 = v_EQ2_0_out0;
assign v_Q0_27_out0 = v__119_out0;
assign v_EQ6_49_out0 = v__14_out1 == 4'h5;
assign v_EQ9_63_out0 = v__14_out1 == 4'h3;
assign v_EQ8_67_out0 = v__14_out1 == 4'h7;
assign v_EQ11_68_out0 = v__14_out1 == 4'h1;
assign v_ADRESS_71_out0 = v__14_out0;
assign v_START_92_out0 = v_EQ4_25_out0;
assign v_EXEC2LS_95_out0 = v_EQ3_192_out0;
assign v_EQ7_105_out0 = v__14_out1 == 4'h6;
assign v_EQ5_118_out0 = v__14_out1 == 4'h4;
assign v_EQ3_136_out0 = v__14_out1 == 4'h2;
assign v_G1_31_out0 = ! v_Q0_27_out0;
assign v_JMI_47_out0 = v_EQ6_49_out0;
assign v_ADRESS_61_out0 = v_ADRESS_71_out0;
assign v_G2_78_out0 = v_EQ9_63_out0 || v_EQ10_59_out0;
assign v_FLOAT_111_out0 = v_EQ3_136_out0;
assign v_G2_121_out0 = ! v_Q1_18_out0;
assign v_EXEC1LS_122_out0 = v_EXEC1LS_22_out0;
assign v_G13_133_out0 = v_Q0_27_out0 && v_Q1_18_out0;
assign v_JMP_143_out0 = v_EQ5_118_out0;
assign v_STP_150_out0 = v_EQ8_67_out0;
assign v_JEQ_153_out0 = v_EQ7_105_out0;
assign v_EXEC2LS_173_out0 = v_EXEC2LS_95_out0;
assign v_G1_177_out0 = v_EQ1_19_out0 || v_EQ9_63_out0;
assign v_START_186_out0 = v_START_92_out0;
assign v_NORMAL_188_out0 = v_NORMAL_13_out0;
assign v_STP_3_out0 = v_STP_150_out0;
assign v_START_20_out0 = v_START_186_out0;
assign v_G7_35_out0 = v_G1_31_out0 && v_Q1_18_out0;
assign v_UART_42_out0 = v_G2_78_out0;
assign v_G3_48_out0 = v_EQ11_68_out0 || v_G1_177_out0;
assign v_JEQ_55_out0 = v_JEQ_153_out0;
assign v_EXEC2LS_99_out0 = v_EXEC2LS_173_out0;
assign v_JMP_100_out0 = v_JMP_143_out0;
assign v_JUMPADRESS_126_out0 = v_ADRESS_61_out0;
assign v_EXEC1_130_out0 = v_EXEC1LS_122_out0;
assign v_FLOAT_138_out0 = v_FLOAT_111_out0;
assign v_NORMAL_144_out0 = v_NORMAL_188_out0;
assign v_EXEC1LS_154_out0 = v_EXEC1LS_122_out0;
assign v_G5_171_out0 = v_Q0_27_out0 && v_G2_121_out0;
assign v_JMI_185_out0 = v_JMI_47_out0;
assign v_G3_194_out0 = v_G1_31_out0 && v_G2_121_out0;
assign v_JMI_9_out0 = v_JMI_185_out0;
assign v_STALL_21_out0 = v_G3_48_out0;
assign v_JMP_24_out0 = v_JMP_100_out0;
assign v_G6_87_out0 = v_G3_194_out0 || v_G7_35_out0;
assign v_G3_89_out0 = v_FLOAT_138_out0 && v_NORMAL_188_out0;
assign v_JMI_97_out0 = v_JMI_185_out0;
assign v_JEQ_109_out0 = v_JEQ_55_out0;
assign v_JUMPADRESS_115_out0 = v_JUMPADRESS_126_out0;
assign v_JMP_132_out0 = v_JMP_100_out0;
assign v_JEQ_142_out0 = v_JEQ_55_out0;
assign v_STP_151_out0 = v_STP_3_out0;
assign v_EXEC1_164_out0 = v_EXEC1_130_out0;
assign v_UART_169_out0 = v_UART_42_out0;
assign v_STP_172_out0 = v_STP_3_out0;
assign v_STALL_39_out0 = v_STALL_21_out0;
assign v_G15_43_out0 = !(v_EXEC1_164_out0 || v_FF1_2_out0);
assign v_G4_117_out0 = v_JEQZ_91_out0 && v_JEQ_142_out0;
assign v_STALL_125_out0 = v_STALL_21_out0;
assign v_G5_157_out0 = v_JMIN_33_out0 && v_JMI_97_out0;
assign v_STP_180_out0 = v_STP_151_out0;
assign v_G9_34_out0 = ! v_STALL_125_out0;
assign v_STALL_145_out0 = v_STALL_39_out0;
assign v_G4_146_out0 = v_G5_171_out0 && v_STALL_125_out0;
assign v_G12_159_out0 = ! v_STP_180_out0;
assign v_G11_189_out0 = v_EXEC1_164_out0 || v_STP_180_out0;
assign v_G2_195_out0 = v_JMP_24_out0 || v_G5_157_out0;
assign v_G8_40_out0 = v_G7_35_out0 || v_G4_146_out0;
assign v_G11_74_out0 = v_G5_171_out0 && v_G9_34_out0;
assign v_SUB_88_out0 = v_G11_189_out0;
assign v_G3_107_out0 = v_G2_195_out0 || v_G4_117_out0;
assign v_G5_15_out0 = ((v__103_out0 && !v_SUB_88_out0) || (!v__103_out0) && v_SUB_88_out0);
assign v_G8_53_out0 = ((v__11_out0 && !v_SUB_88_out0) || (!v__11_out0) && v_SUB_88_out0);
assign v_JUMP_54_out0 = v_G3_107_out0;
assign v_G9_60_out0 = ((v__56_out0 && !v_SUB_88_out0) || (!v__56_out0) && v_SUB_88_out0);
assign v_G6_65_out0 = ((v__52_out0 && !v_SUB_88_out0) || (!v__52_out0) && v_SUB_88_out0);
assign v_G11_72_out0 = ((v__4_out0 && !v_SUB_88_out0) || (!v__4_out0) && v_SUB_88_out0);
assign v_G3_73_out0 = ((v__17_out0 && !v_SUB_88_out0) || (!v__17_out0) && v_SUB_88_out0);
assign v_G10_76_out0 = ((v__181_out0 && !v_SUB_88_out0) || (!v__181_out0) && v_SUB_88_out0);
assign v_G2_101_out0 = ((v__93_out0 && !v_SUB_88_out0) || (!v__93_out0) && v_SUB_88_out0);
assign v_G12_113_out0 = ((v__45_out0 && !v_SUB_88_out0) || (!v__45_out0) && v_SUB_88_out0);
assign v_G7_116_out0 = ((v__187_out0 && !v_SUB_88_out0) || (!v__187_out0) && v_SUB_88_out0);
assign v_G12_147_out0 = v_G11_74_out0 && v_G2_121_out0;
assign v_G1_152_out0 = ((v__193_out0 && !v_SUB_88_out0) || (!v__193_out0) && v_SUB_88_out0);
assign v_G4_183_out0 = ((v__12_out0 && !v_SUB_88_out0) || (!v__12_out0) && v_SUB_88_out0);
assign v_G14_32_out0 = v_G15_43_out0 && v_JUMP_54_out0;
assign v__36_out0 = { v_G1_152_out0,v_G2_101_out0 };
assign v_G10_38_out0 = v_G6_87_out0 || v_G12_147_out0;
assign v__62_out0 = { v__36_out0,v_G3_73_out0 };
assign v_MUX1_165_out0 = v_G14_32_out0 ? v_JUMPADRESS_115_out0 : v_REG1_23_out0;
assign v_G14_184_out0 = v_G10_38_out0 || v_G13_133_out0;
assign v__90_out0 = { v__62_out0,v_G4_183_out0 };
assign v__175_out0 = { v_G14_184_out0,v_G8_40_out0 };
assign v_D_26_out0 = v__175_out0;
assign v__120_out0 = { v__90_out0,v_G5_15_out0 };
assign v__10_out0 = { v__120_out0,v_G6_65_out0 };
assign v__112_out0 = v_D_26_out0[0:0];
assign v__112_out1 = v_D_26_out0[1:1];
assign v__7_out0 = { v__10_out0,v_G7_116_out0 };
assign v__140_out0 = { v__7_out0,v_G8_53_out0 };
assign v__84_out0 = { v__140_out0,v_G9_60_out0 };
assign v__77_out0 = { v__84_out0,v_G10_76_out0 };
assign v__114_out0 = { v__77_out0,v_G11_72_out0 };
assign v__166_out0 = { v__114_out0,v_G12_113_out0 };
assign v_ADDER_IN_174_out0 = v__166_out0;
assign {v_A1_128_out1,v_A1_128_out0 } = v_MUX1_165_out0 + v_ADDER_IN_174_out0 + v_G11_189_out0;
assign v_COUT_6_out0 = v_A1_128_out1;
assign v_MUX4_79_out0 = v_BYTE_READY_85_out0 ? v_C1_66_out0 : v_A1_128_out0;
assign v_MUX3_149_out0 = v_STP_180_out0 ? v_A1_128_out0 : v_MUX1_165_out0;
assign v_PC_COUNTER_NEXT_131_out0 = v_MUX3_149_out0;
assign v_PC_COUNTER_1_out0 = v_PC_COUNTER_NEXT_131_out0;
assign v_MUX1_64_out0 = v_EXEC1LS_122_out0 ? v_RAMADDRESSMUX_123_out0 : v_PC_COUNTER_NEXT_131_out0;
assign v_MUX3_98_out0 = v_BYTE_READY_129_out0 ? v_C2_163_out0 : v_MUX1_64_out0;
assign v__141_out0 = { v_PC_COUNTER_1_out0,v_C1_50_out0 };
assign v_MUX2_96_out0 = v_BYTE_READY_129_out0 ? v__141_out0 : v_RAM_IN_16_out0;
assign v_NEXTADD_156_out0 = v_MUX3_98_out0;


endmodule



    module v_ROM1_225(q, a, clk);
    output reg [0:0] q;
    input [11:0] a;
    reg [0:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end
    begin
        rom[0] = 0;
rom[1] = 1;
rom[2] = 0;
rom[3] = 0;
rom[4] = 0;
rom[5] = 0;
rom[6] = 0;
rom[7] = 0;
rom[8] = 0;
rom[9] = 1;
rom[10] = 1;
rom[11] = 1;
rom[12] = 0;
rom[13] = 0;
rom[14] = 1;
rom[15] = 0;
rom[16] = 0;
rom[17] = 0;
rom[18] = 0;
rom[19] = 0;
rom[20] = 0;
rom[21] = 1;
rom[22] = 1;
rom[23] = 1;
rom[24] = 1;
rom[25] = 0;
rom[26] = 0;
rom[27] = 0;
rom[28] = 0;
rom[29] = 0;
rom[30] = 0;
rom[31] = 1;
rom[32] = 1;
rom[33] = 1;
rom[34] = 1;
rom[35] = 1;
rom[36] = 1;
rom[37] = 1;
rom[38] = 1;
rom[39] = 1;
rom[40] = 1;
rom[41] = 1;
rom[42] = 1;
rom[43] = 1;
rom[44] = 1;
rom[45] = 1;
rom[46] = 1;
rom[47] = 1;
rom[48] = 1;
rom[49] = 1;
rom[50] = 1;
rom[51] = 1;
rom[52] = 1;
rom[53] = 1;
rom[54] = 1;
rom[55] = 1;
rom[56] = 1;
rom[57] = 1;
rom[58] = 1;
rom[59] = 1;
rom[60] = 1;
rom[61] = 1;
rom[62] = 1;
rom[63] = 1;
rom[64] = 1;
rom[65] = 1;
rom[66] = 1;
rom[67] = 1;
rom[68] = 1;
rom[69] = 1;
rom[70] = 1;
rom[71] = 1;
rom[72] = 1;
rom[73] = 1;
rom[74] = 1;
rom[75] = 1;
rom[76] = 1;
rom[77] = 1;
rom[78] = 1;
rom[79] = 1;
rom[80] = 1;
rom[81] = 1;
rom[82] = 1;
rom[83] = 1;
rom[84] = 1;
rom[85] = 1;
rom[86] = 1;
rom[87] = 1;
rom[88] = 1;
rom[89] = 1;
rom[90] = 1;
rom[91] = 1;
rom[92] = 1;
rom[93] = 1;
rom[94] = 1;
rom[95] = 1;
    end
     

    module v_RAM1_930(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 724;
ram[1] = 1753;
ram[2] = 2782;
ram[3] = 3811;
ram[4] = 16393;
ram[5] = 15360;
ram[6] = 12629;
ram[7] = 8260;
ram[8] = 2624;
ram[9] = 8192;
ram[10] = 36865;
ram[11] = 32770;
ram[12] = 36867;
ram[13] = 0;
ram[14] = 0;
ram[15] = 0;
ram[16] = 0;
ram[17] = 49668;
ram[18] = 52738;
ram[19] = 35840;
ram[20] = 3585;
ram[21] = 3074;
ram[22] = 3288;
ram[32] = 12801;
ram[33] = 35840;
ram[34] = 15362;
ram[35] = 3280;
ram[37] = 1792;
ram[127] = 49775;
ram[255] = 1058;
ram[256] = 32768;
ram[257] = 61440;
ram[258] = 258;
ram[2038] = 198;
ram[2039] = 3274;
ram[2040] = 12801;
ram[2041] = 3790;
ram[2042] = 35840;
ram[2043] = 15362;
ram[2044] = 3278;
ram[2045] = 710;
ram[2046] = 3786;
    end
    endmodule

    
module main (
	clk,
	v_DIV_INST_1133_out0,
	v_TX_OVERFLOW_1184_out0,
	v_RECEIVE_REGISTER_2841_out0,
	v_RD_1006_out0,
	v_STP_6646_out0,
	v_MULTI_OPCODE_3499_out0,
	v_RM_1555_out0,
	v_WEN_MULTI_2240_out0,
	v_BYTE_READY_RX_6654_out0,
	v_TRANSMISSION_DATA_1422_out0,
	v_INSTRCUTION_1926_out0,
	v_TRANSMITER_1BIT_1296_out0,
	v_MULTI_OUT_1589_out0);
input clk;
input v_DIV_INST_1133_out0;
output  [15:0] v_MULTI_OUT_1589_out0;
output  [15:0] v_RM_1555_out0;
output  [1:0] v_RD_1006_out0;
output  [7:0] v_RECEIVE_REGISTER_2841_out0;
output  [7:0] v_TRANSMISSION_DATA_1422_out0;
output v_BYTE_READY_RX_6654_out0;
output v_INSTRCUTION_1926_out0;
output v_MULTI_OPCODE_3499_out0;
output v_STP_6646_out0;
output v_TRANSMITER_1BIT_1296_out0;
output v_TX_OVERFLOW_1184_out0;
output v_WEN_MULTI_2240_out0;
reg  [11:0] v_REG1_210_out0 = 12'h0;
reg  [11:0] v_REG1_3500_out0 = 12'h0;
reg  [15:0] v_IHOLD_REGISTER_983_out0 = 16'h0;
reg  [15:0] v_REG0_5368_out0 = 16'h0;
reg  [15:0] v_REG1_1128_out0 = 16'h0;
reg  [15:0] v_REG1_6571_out0 = 16'h0;
reg  [15:0] v_REG2_6035_out0 = 16'h0;
reg  [15:0] v_REG3_2317_out0 = 16'h0;
reg  [1:0] v_REG1_5108_out0 = 2'h0;
reg  [7:0] v_REG1_1306_out0 = 8'h0;
reg  [7:0] v_REG1_5190_out0 = 8'h0;
reg v_FF1_2303_out0 = 1'b0;
reg v_FF1_2304_out0 = 1'b0;
reg v_FF1_2305_out0 = 1'b0;
reg v_FF1_2306_out0 = 1'b0;
reg v_FF1_2307_out0 = 1'b0;
reg v_FF1_2308_out0 = 1'b0;
reg v_FF1_2309_out0 = 1'b0;
reg v_FF1_2310_out0 = 1'b0;
reg v_FF1_26_out0 = 1'b0;
reg v_FF1_5090_out0 = 1'b0;
reg v_FF1_5442_out0 = 1'b0;
reg v_FF1_6658_out0 = 1'b0;
reg v_FF1_956_out0 = 1'b0;
reg v_FF2_1362_out0 = 1'b0;
reg v_FF2_1383_out0 = 1'b0;
reg v_FF2_43_out0 = 1'b0;
reg v_FF2_5444_out0 = 1'b0;
reg v_FF3_5175_out0 = 1'b0;
reg v_FF3_5435_out0 = 1'b0;
reg v_FF4_226_out0 = 1'b0;
reg v_FF5_3484_out0 = 1'b0;
reg v_FF6_58_out0 = 1'b0;
reg v_FF7_1302_out0 = 1'b0;
reg v_FF7_1303_out0 = 1'b0;
reg v_FF7_2334_out0 = 1'b0;
reg v_FF8_5337_out0 = 1'b0;
reg v_FF8_5338_out0 = 1'b0;
reg v_FF8_5523_out0 = 1'b0;
reg v_FF9_4333_out0 = 1'b0;
reg v_REG1_5479_out0 = 1'b0;
wire  [10:0] v_C1_294_out0;
wire  [10:0] v_IN1_1067_out0;
wire  [10:0] v_IN1_1391_out0;
wire  [10:0] v_IN1_5410_out0;
wire  [10:0] v_IN1_6754_out0;
wire  [10:0] v_IN_6733_out0;
wire  [10:0] v_MUX1_1171_out0;
wire  [10:0] v_MUX1_3504_out0;
wire  [10:0] v_MUX1_3784_out0;
wire  [10:0] v_MUX2_95_out0;
wire  [10:0] v_MUX3_6560_out0;
wire  [10:0] v_MUX4_271_out0;
wire  [10:0] v_MUX5_6734_out0;
wire  [10:0] v_OP2_SIG11_2357_out0;
wire  [10:0] v_OP2_SIG11_8_out0;
wire  [10:0] v_OP2_SIG_6561_out0;
wire  [10:0] v_OP2_SIG_NEW_5507_out0;
wire  [10:0] v_OP2_SIG_NEW_5520_out0;
wire  [10:0] v_OUT1_1601_out0;
wire  [10:0] v_OUT1_1878_out0;
wire  [10:0] v_OUT1_916_out0;
wire  [10:0] v_OUT1_964_out0;
wire  [10:0] v_Q_5096_out0;
wire  [10:0] v_Q_5097_out0;
wire  [10:0] v_RD_SIG11_3498_out0;
wire  [10:0] v_RD_SIG11_4356_out0;
wire  [10:0] v_RD_SIG_56_out0;
wire  [10:0] v_RD_SIG_NEW_4310_out0;
wire  [10:0] v_RD_SIG_NEW_5348_out0;
wire  [10:0] v_SEL2_6650_out0;
wire  [10:0] v_SHIFTED_SIG_5314_out0;
wire  [10:0] v_SHIFTED_SIG_6716_out0;
wire  [10:0] v_SIG_RD_11bit_1605_out0;
wire  [10:0] v_SIG_RM_11bit_3384_out0;
wire  [10:0] v_SIG_TO_SHIFT_2861_out0;
wire  [10:0] v_SIG_TO_SHIFT_5273_out0;
wire  [10:0] v__1000_out0;
wire  [10:0] v__1001_out0;
wire  [10:0] v__1002_out0;
wire  [10:0] v__1068_out0;
wire  [10:0] v__1352_out0;
wire  [10:0] v__1384_out0;
wire  [10:0] v__1385_out0;
wire  [10:0] v__1450_out0;
wire  [10:0] v__2242_out0;
wire  [10:0] v__2311_out0;
wire  [10:0] v__3790_out0;
wire  [10:0] v__6559_out0;
wire  [10:0] v__6642_out0;
wire  [10:0] v__6778_out0;
wire  [10:0] v__988_out0;
wire  [10:0] v__989_out0;
wire  [10:0] v__990_out0;
wire  [10:0] v__991_out0;
wire  [10:0] v__992_out0;
wire  [10:0] v__993_out0;
wire  [10:0] v__994_out0;
wire  [10:0] v__995_out0;
wire  [10:0] v__996_out0;
wire  [10:0] v__997_out0;
wire  [10:0] v__998_out0;
wire  [10:0] v__999_out0;
wire  [10:0] v_shifted1_1300_out0;
wire  [11:0] v_A1_3446_out0;
wire  [11:0] v_A1_5433_out0;
wire  [11:0] v_ADDER_IN_5411_out0;
wire  [11:0] v_ADRESS_1141_out0;
wire  [11:0] v_ADRESS_1239_out0;
wire  [11:0] v_A_5323_out0;
wire  [11:0] v_C1_1182_out0;
wire  [11:0] v_C1_1564_out0;
wire  [11:0] v_C2_1176_out0;
wire  [11:0] v_C2_5297_out0;
wire  [11:0] v_C_883_out0;
wire  [11:0] v_EA_6661_out0;
wire  [11:0] v_JUMPADRESS_2316_out0;
wire  [11:0] v_JUMPADRESS_3419_out0;
wire  [11:0] v_MULTI_PRODUCT_3485_out0;
wire  [11:0] v_MUX1_1169_out0;
wire  [11:0] v_MUX1_5302_out0;
wire  [11:0] v_MUX2_6726_out0;
wire  [11:0] v_MUX3_1571_out0;
wire  [11:0] v_MUX3_5092_out0;
wire  [11:0] v_MUX4_1295_out0;
wire  [11:0] v_MUX8_6790_out0;
wire  [11:0] v_NEXTADD_5180_out0;
wire  [11:0] v_NEXTADRESS_882_out0;
wire  [11:0] v_NOUSED_6647_out0;
wire  [11:0] v_PC_COUNTER_16_out0;
wire  [11:0] v_PC_COUNTER_NEXT_3468_out0;
wire  [11:0] v_RAMADDRESSMUX_3375_out0;
wire  [11:0] v_RAMADDRMUX_1088_out0;
wire  [11:0] v_RAMADDRMUX_48_out0;
wire  [11:0] v_RAMADDRMUX_5187_out0;
wire  [11:0] v_RAM_ADDRESS_MUX_4332_out0;
wire  [11:0] v_SEL7_2367_out0;
wire  [11:0] v_SEL8_5260_out0;
wire  [11:0] v__112_out0;
wire  [11:0] v__1175_out0;
wire  [11:0] v__1187_out0;
wire  [11:0] v__1364_out0;
wire  [11:0] v__1365_out0;
wire  [11:0] v__1366_out0;
wire  [11:0] v__1367_out0;
wire  [11:0] v__1368_out0;
wire  [11:0] v__1369_out0;
wire  [11:0] v__1370_out0;
wire  [11:0] v__1371_out0;
wire  [11:0] v__1372_out0;
wire  [11:0] v__1373_out0;
wire  [11:0] v__1374_out0;
wire  [11:0] v__1375_out0;
wire  [11:0] v__1376_out0;
wire  [11:0] v__1377_out0;
wire  [11:0] v__1378_out0;
wire  [11:0] v__1479_out0;
wire  [11:0] v__2193_out1;
wire  [11:0] v__2237_out1;
wire  [11:0] v__2865_out0;
wire  [11:0] v__3490_out0;
wire  [11:0] v__5307_out0;
wire  [11:0] v__5482_out0;
wire  [11:0] v__5483_out0;
wire  [11:0] v__55_out0;
wire  [11:0] v__6554_out1;
wire  [12:0] v__1557_out0;
wire  [12:0] v__1558_out0;
wire  [12:0] v__2867_out0;
wire  [12:0] v__4830_out0;
wire  [12:0] v__84_out0;
wire  [12:0] v__891_out0;
wire  [12:0] v__892_out0;
wire  [12:0] v__893_out0;
wire  [12:0] v__894_out0;
wire  [12:0] v__895_out0;
wire  [12:0] v__896_out0;
wire  [12:0] v__897_out0;
wire  [12:0] v__898_out0;
wire  [12:0] v__899_out0;
wire  [12:0] v__900_out0;
wire  [12:0] v__901_out0;
wire  [12:0] v__902_out0;
wire  [12:0] v__903_out0;
wire  [12:0] v__904_out0;
wire  [12:0] v__905_out0;
wire  [13:0] v__2190_out1;
wire  [13:0] v__2220_out0;
wire  [13:0] v__2221_out0;
wire  [13:0] v__2222_out0;
wire  [13:0] v__2223_out0;
wire  [13:0] v__2224_out0;
wire  [13:0] v__2225_out0;
wire  [13:0] v__2226_out0;
wire  [13:0] v__2227_out0;
wire  [13:0] v__2228_out0;
wire  [13:0] v__2229_out0;
wire  [13:0] v__2230_out0;
wire  [13:0] v__2231_out0;
wire  [13:0] v__2232_out0;
wire  [13:0] v__2233_out0;
wire  [13:0] v__2234_out0;
wire  [13:0] v__2352_out1;
wire  [13:0] v__264_out0;
wire  [13:0] v__304_out1;
wire  [13:0] v__5300_out0;
wire  [13:0] v__5437_out0;
wire  [13:0] v__5440_out0;
wire  [13:0] v__89_out0;
wire  [13:0] v__90_out0;
wire  [14:0] v_CIN_1148_out0;
wire  [14:0] v_REST_83_out0;
wire  [14:0] v__1084_out0;
wire  [14:0] v__1407_out1;
wire  [14:0] v__1456_out1;
wire  [14:0] v__2358_out0;
wire  [14:0] v__2370_out1;
wire  [14:0] v__5102_out0;
wire  [14:0] v__5149_out0;
wire  [14:0] v__5150_out0;
wire  [14:0] v__5243_out0;
wire  [14:0] v__5244_out0;
wire  [14:0] v__5245_out0;
wire  [14:0] v__5246_out0;
wire  [14:0] v__5247_out0;
wire  [14:0] v__5248_out0;
wire  [14:0] v__5249_out0;
wire  [14:0] v__5250_out0;
wire  [14:0] v__5251_out0;
wire  [14:0] v__5252_out0;
wire  [14:0] v__5253_out0;
wire  [14:0] v__5254_out0;
wire  [14:0] v__5255_out0;
wire  [14:0] v__5256_out0;
wire  [14:0] v__5257_out0;
wire  [14:0] v__5367_out1;
wire  [14:0] v__5528_out0;
wire  [14:0] v__5559_out0;
wire  [14:0] v__6753_out0;
wire  [15:0] v_16BIT_WORD_ANSWER_4340_out0;
wire  [15:0] v_A1_1547_out0;
wire  [15:0] v_A1_1879_out0;
wire  [15:0] v_A4_5526_out0;
wire  [15:0] v_A5_929_out0;
wire  [15:0] v_A6_5152_out0;
wire  [15:0] v_A8_5490_out0;
wire  [15:0] v_ADDER_IN_4303_out0;
wire  [15:0] v_ADDER_IN_4304_out0;
wire  [15:0] v_ALUOUT_2195_out0;
wire  [15:0] v_ALUOUT_2249_out0;
wire  [15:0] v_ALUOUT_4357_out0;
wire  [15:0] v_ALUOUT_5181_out0;
wire  [15:0] v_ALUOUT_5439_out0;
wire  [15:0] v_ANDOUT_305_out0;
wire  [15:0] v_ANDOUT_306_out0;
wire  [15:0] v_A_5066_out0;
wire  [15:0] v_A_5067_out0;
wire  [15:0] v_A_5537_out0;
wire  [15:0] v_A_5538_out0;
wire  [15:0] v_B_1629_out0;
wire  [15:0] v_C11_2218_out0;
wire  [15:0] v_C13_1065_out0;
wire  [15:0] v_C15_847_out0;
wire  [15:0] v_C5_1312_out0;
wire  [15:0] v_C7_912_out0;
wire  [15:0] v_CIN_1147_out0;
wire  [15:0] v_CIN_1149_out0;
wire  [15:0] v_CIN_1150_out0;
wire  [15:0] v_CIN_1151_out0;
wire  [15:0] v_CIN_1152_out0;
wire  [15:0] v_CIN_1153_out0;
wire  [15:0] v_CIN_1154_out0;
wire  [15:0] v_CIN_1155_out0;
wire  [15:0] v_CIN_1156_out0;
wire  [15:0] v_CIN_1157_out0;
wire  [15:0] v_CIN_1158_out0;
wire  [15:0] v_CIN_1159_out0;
wire  [15:0] v_CIN_1160_out0;
wire  [15:0] v_CIN_1161_out0;
wire  [15:0] v_COUT_5371_out0;
wire  [15:0] v_COUT_5372_out0;
wire  [15:0] v_COUT_5373_out0;
wire  [15:0] v_COUT_5374_out0;
wire  [15:0] v_COUT_5375_out0;
wire  [15:0] v_COUT_5376_out0;
wire  [15:0] v_COUT_5377_out0;
wire  [15:0] v_COUT_5378_out0;
wire  [15:0] v_COUT_5379_out0;
wire  [15:0] v_COUT_5380_out0;
wire  [15:0] v_COUT_5381_out0;
wire  [15:0] v_COUT_5382_out0;
wire  [15:0] v_COUT_5383_out0;
wire  [15:0] v_COUT_5384_out0;
wire  [15:0] v_COUT_5385_out0;
wire  [15:0] v_DIN3_5083_out0;
wire  [15:0] v_DIN_1105_out0;
wire  [15:0] v_DIN_4828_out0;
wire  [15:0] v_DOUT1_591_out0;
wire  [15:0] v_DOUT2_848_out0;
wire  [15:0] v_FLOATING_REGISTER_IN_275_out0;
wire  [15:0] v_IN_1145_out0;
wire  [15:0] v_IN_1299_out0;
wire  [15:0] v_IN_2840_out0;
wire  [15:0] v_IN_332_out0;
wire  [15:0] v_IN_4348_out0;
wire  [15:0] v_IN_5124_out0;
wire  [15:0] v_IN_51_out0;
wire  [15:0] v_IN_5542_out0;
wire  [15:0] v_IN_6557_out0;
wire  [15:0] v_IN_6677_out0;
wire  [15:0] v_IN_6792_out0;
wire  [15:0] v_IN_960_out0;
wire  [15:0] v_IN_96_out0;
wire  [15:0] v_IR_1380_out0;
wire  [15:0] v_IR_1413_out0;
wire  [15:0] v_IR_3489_out0;
wire  [15:0] v_IR_5321_out0;
wire  [15:0] v_IR_54_out0;
wire  [15:0] v_IR_6640_out0;
wire  [15:0] v_IR_915_out0;
wire  [15:0] v_KEXTEND_6567_out0;
wire  [15:0] v_LS_REGIN_1606_out0;
wire  [15:0] v_MULTI_OUT_6706_out0;
wire  [15:0] v_MULTI_REGIN_1399_out0;
wire  [15:0] v_MUX11_6771_out0;
wire  [15:0] v_MUX12_840_out0;
wire  [15:0] v_MUX1_1235_out0;
wire  [15:0] v_MUX1_1326_out0;
wire  [15:0] v_MUX1_19_out0;
wire  [15:0] v_MUX1_2364_out0;
wire  [15:0] v_MUX1_3_out0;
wire  [15:0] v_MUX1_4337_out0;
wire  [15:0] v_MUX1_5143_out0;
wire  [15:0] v_MUX1_5484_out0;
wire  [15:0] v_MUX1_849_out0;
wire  [15:0] v_MUX1_921_out0;
wire  [15:0] v_MUX2_1140_out0;
wire  [15:0] v_MUX2_1561_out0;
wire  [15:0] v_MUX2_1585_out0;
wire  [15:0] v_MUX2_2252_out0;
wire  [15:0] v_MUX2_5334_out0;
wire  [15:0] v_MUX2_579_out0;
wire  [15:0] v_MUX2_588_out0;
wire  [15:0] v_MUX2_6563_out0;
wire  [15:0] v_MUX3_1004_out0;
wire  [15:0] v_MUX3_1483_out0;
wire  [15:0] v_MUX3_1527_out0;
wire  [15:0] v_MUX3_155_out0;
wire  [15:0] v_MUX3_3371_out0;
wire  [15:0] v_MUX3_3474_out0;
wire  [15:0] v_MUX3_4267_out0;
wire  [15:0] v_MUX3_6570_out0;
wire  [15:0] v_MUX4_1087_out0;
wire  [15:0] v_MUX4_186_out0;
wire  [15:0] v_MUX4_3448_out0;
wire  [15:0] v_MUX4_5179_out0;
wire  [15:0] v_MUX4_6651_out0;
wire  [15:0] v_MUX4_6_out0;
wire  [15:0] v_MUX5_1265_out0;
wire  [15:0] v_MUX5_1270_out0;
wire  [15:0] v_MUX5_1607_out0;
wire  [15:0] v_MUX5_3445_out0;
wire  [15:0] v_MUX5_4349_out0;
wire  [15:0] v_MUX5_5220_out0;
wire  [15:0] v_MUX5_581_out0;
wire  [15:0] v_MUX6_1142_out0;
wire  [15:0] v_MUX7_572_out0;
wire  [15:0] v_MUX8_932_out0;
wire  [15:0] v_M_REGIN_135_out0;
wire  [15:0] v_OP1_1005_out0;
wire  [15:0] v_OP1_1454_out0;
wire  [15:0] v_OP1_1900_out0;
wire  [15:0] v_OP2_1132_out0;
wire  [15:0] v_OP2_1397_out0;
wire  [15:0] v_OP2_1921_out0;
wire  [15:0] v_OP2_5292_out0;
wire  [15:0] v_OP2_5489_out0;
wire  [15:0] v_OUT_1146_out0;
wire  [15:0] v_OUT_1394_out0;
wire  [15:0] v_OUT_224_out0;
wire  [15:0] v_OUT_3787_out0;
wire  [15:0] v_OUT_3788_out0;
wire  [15:0] v_OUT_4355_out0;
wire  [15:0] v_OUT_5062_out0;
wire  [15:0] v_OUT_5529_out0;
wire  [15:0] v_OUT_557_out0;
wire  [15:0] v_OUT_6029_out0;
wire  [15:0] v_R0TEST_1552_out0;
wire  [15:0] v_R0TEST_3439_out0;
wire  [15:0] v_R0_1237_out0;
wire  [15:0] v_R0_1392_out0;
wire  [15:0] v_R0_828_out0;
wire  [15:0] v_R1TEST_5162_out0;
wire  [15:0] v_R1TEST_5168_out0;
wire  [15:0] v_R1_1003_out0;
wire  [15:0] v_R1_1282_out0;
wire  [15:0] v_R1_4311_out0;
wire  [15:0] v_R2TEST_5270_out0;
wire  [15:0] v_R2TEST_5407_out0;
wire  [15:0] v_R2_1484_out0;
wire  [15:0] v_R2_5194_out0;
wire  [15:0] v_R2_5364_out0;
wire  [15:0] v_R3TEST_1400_out0;
wire  [15:0] v_R3TEST_61_out0;
wire  [15:0] v_R3_20_out0;
wire  [15:0] v_R3_2273_out0;
wire  [15:0] v_R3_38_out0;
wire  [15:0] v_RAM1_930_out0;
wire  [15:0] v_RAMDOUT_1177_out0;
wire  [15:0] v_RAMDOUT_1478_out0;
wire  [15:0] v_RAMDOUT_14_out0;
wire  [15:0] v_RAM_IN_116_out0;
wire  [15:0] v_RAM_OUT_200_out0;
wire  [15:0] v_RAM_OUT_3506_out0;
wire  [15:0] v_RAM_OUT_5519_out0;
wire  [15:0] v_RAM_OUT_5521_out0;
wire  [15:0] v_RAM_OUT_855_out0;
wire  [15:0] v_RDOUT_1360_out0;
wire  [15:0] v_RD_1896_out0;
wire  [15:0] v_RD_2362_out0;
wire  [15:0] v_RD_245_out0;
wire  [15:0] v_RD_297_out0;
wire  [15:0] v_RD_FLOATING_1379_out0;
wire  [15:0] v_RD_MULTI_25_out0;
wire  [15:0] v_REGDIN_5432_out0;
wire  [15:0] v_REGISTER_INPUT_6543_out0;
wire  [15:0] v_REGISTER_OUTPUT_6728_out0;
wire  [15:0] v_REGISTER_OUT_5064_out0;
wire  [15:0] v_RMN_6619_out0;
wire  [15:0] v_RM_1420_out0;
wire  [15:0] v_RM_1591_out0;
wire  [15:0] v_RM_2217_out0;
wire  [15:0] v_RM_4298_out0;
wire  [15:0] v_RM_5445_out0;
wire  [15:0] v_RM_5446_out0;
wire  [15:0] v_RM_5447_out0;
wire  [15:0] v_RM_5448_out0;
wire  [15:0] v_RM_5449_out0;
wire  [15:0] v_RM_5450_out0;
wire  [15:0] v_RM_5451_out0;
wire  [15:0] v_RM_5452_out0;
wire  [15:0] v_RM_5453_out0;
wire  [15:0] v_RM_5454_out0;
wire  [15:0] v_RM_5455_out0;
wire  [15:0] v_RM_5456_out0;
wire  [15:0] v_RM_5457_out0;
wire  [15:0] v_RM_5458_out0;
wire  [15:0] v_RM_5459_out0;
wire  [15:0] v_RM_5496_out0;
wire  [15:0] v_RM_6657_out0;
wire  [15:0] v_RM_6701_out0;
wire  [15:0] v_RM_6773_out0;
wire  [15:0] v_RM_MULTI_105_out0;
wire  [15:0] v_RM_MULTI_313_out0;
wire  [15:0] v_SUM1_6516_out0;
wire  [15:0] v_XOR1_5534_out0;
wire  [15:0] v_XOR2_2192_out0;
wire  [15:0] v_XOR3_6702_out0;
wire  [15:0] v__1307_out0;
wire  [15:0] v__1363_out0;
wire  [15:0] v__1549_out0;
wire  [15:0] v__165_out0;
wire  [15:0] v__195_out0;
wire  [15:0] v__2276_out0;
wire  [15:0] v__2299_out0;
wire  [15:0] v__3374_out0;
wire  [15:0] v__3476_out0;
wire  [15:0] v__3492_out0;
wire  [15:0] v__3494_out0;
wire  [15:0] v__3523_out0;
wire  [15:0] v__3753_out0;
wire  [15:0] v__3754_out0;
wire  [15:0] v__4281_out0;
wire  [15:0] v__4824_out0;
wire  [15:0] v__5094_out0;
wire  [15:0] v__5146_out0;
wire  [15:0] v__5170_out0;
wire  [15:0] v__5320_out0;
wire  [15:0] v__5386_out0;
wire  [15:0] v__5387_out0;
wire  [15:0] v__5388_out0;
wire  [15:0] v__5389_out0;
wire  [15:0] v__5390_out0;
wire  [15:0] v__5391_out0;
wire  [15:0] v__5392_out0;
wire  [15:0] v__5393_out0;
wire  [15:0] v__5394_out0;
wire  [15:0] v__5395_out0;
wire  [15:0] v__5396_out0;
wire  [15:0] v__5397_out0;
wire  [15:0] v__5398_out0;
wire  [15:0] v__5399_out0;
wire  [15:0] v__5400_out0;
wire  [15:0] v__5527_out0;
wire  [15:0] v__575_out0;
wire  [15:0] v__592_out0;
wire  [15:0] v__593_out0;
wire  [15:0] v__594_out0;
wire  [15:0] v__64_out0;
wire  [15:0] v__6546_out0;
wire  [15:0] v__6641_out0;
wire  [15:0] v__86_out0;
wire  [15:0] v__913_out0;
wire  [15:0] v__914_out0;
wire  [1:0] v_4BITCOUNTERTRANSIMITER_5539_out0;
wire  [1:0] v_4BITCOUNTER_1419_out0;
wire  [1:0] v_4BITCOUNTER_157_out0;
wire  [1:0] v_4BITCOUNTER_158_out0;
wire  [1:0] v_4BITCOUNTER_2360_out0;
wire  [1:0] v_4BITCOUNTER_4_out0;
wire  [1:0] v_AD1_6785_out0;
wire  [1:0] v_AD2_5266_out0;
wire  [1:0] v_AD3_4269_out0;
wire  [1:0] v_AD3_5161_out0;
wire  [1:0] v_AD3_6545_out0;
wire  [1:0] v_C1_1562_out0;
wire  [1:0] v_C1_3337_out0;
wire  [1:0] v_C1_5558_out0;
wire  [1:0] v_D_1027_out0;
wire  [1:0] v_D_302_out0;
wire  [1:0] v_D_4307_out0;
wire  [1:0] v_MUX1_262_out0;
wire  [1:0] v_MUX2_562_out0;
wire  [1:0] v_M_2295_out0;
wire  [1:0] v_M_3522_out0;
wire  [1:0] v_NOTUSED_1262_out0;
wire  [1:0] v_NOTUSED_217_out0;
wire  [1:0] v_NOTUSED_218_out0;
wire  [1:0] v_Q_5226_out0;
wire  [1:0] v_Q_566_out0;
wire  [1:0] v_ROR_34_out0;
wire  [1:0] v_SHIFT_4263_out0;
wire  [1:0] v_SHIFT_5225_out0;
wire  [1:0] v_SR_184_out0;
wire  [1:0] v_SR_266_out0;
wire  [1:0] v_SR_5221_out0;
wire  [1:0] v_SR_957_out0;
wire  [1:0] v_UARTCOUNTER_1137_out0;
wire  [1:0] v_UART_COUNTER_5328_out0;
wire  [1:0] v_UNUSED_5533_out0;
wire  [1:0] v__1267_out0;
wire  [1:0] v__1406_out0;
wire  [1:0] v__1437_out0;
wire  [1:0] v__1438_out0;
wire  [1:0] v__1566_out0;
wire  [1:0] v__1567_out0;
wire  [1:0] v__1570_out0;
wire  [1:0] v__1594_out0;
wire  [1:0] v__1595_out0;
wire  [1:0] v__188_out0;
wire  [1:0] v__189_out0;
wire  [1:0] v__193_out0;
wire  [1:0] v__194_out0;
wire  [1:0] v__2190_out0;
wire  [1:0] v__2335_out0;
wire  [1:0] v__2336_out0;
wire  [1:0] v__2337_out0;
wire  [1:0] v__2338_out0;
wire  [1:0] v__2339_out0;
wire  [1:0] v__2340_out0;
wire  [1:0] v__2341_out0;
wire  [1:0] v__2342_out0;
wire  [1:0] v__2343_out0;
wire  [1:0] v__2344_out0;
wire  [1:0] v__2345_out0;
wire  [1:0] v__2346_out0;
wire  [1:0] v__2347_out0;
wire  [1:0] v__2348_out0;
wire  [1:0] v__2349_out0;
wire  [1:0] v__2352_out0;
wire  [1:0] v__261_out0;
wire  [1:0] v__304_out0;
wire  [1:0] v__3501_out0;
wire  [1:0] v__3502_out0;
wire  [1:0] v__3525_out0;
wire  [1:0] v__3526_out0;
wire  [1:0] v__5073_out0;
wire  [1:0] v__5074_out0;
wire  [1:0] v__5310_out0;
wire  [1:0] v__5437_out1;
wire  [1:0] v__5441_out0;
wire  [1:0] v__5494_out0;
wire  [1:0] v__559_out0;
wire  [1:0] v__6538_out0;
wire  [1:0] v__6539_out0;
wire  [1:0] v__6678_out0;
wire  [1:0] v__6783_out0;
wire  [1:0] v__6784_out0;
wire  [1:0] v__836_out0;
wire  [1:0] v__954_out0;
wire  [1:0] v__955_out0;
wire  [2:0] v_OP_301_out0;
wire  [2:0] v_OP_5524_out0;
wire  [2:0] v__1163_out0;
wire  [2:0] v__1244_out0;
wire  [2:0] v__1245_out0;
wire  [2:0] v__1246_out0;
wire  [2:0] v__1247_out0;
wire  [2:0] v__1248_out0;
wire  [2:0] v__1249_out0;
wire  [2:0] v__1250_out0;
wire  [2:0] v__1251_out0;
wire  [2:0] v__1252_out0;
wire  [2:0] v__1253_out0;
wire  [2:0] v__1254_out0;
wire  [2:0] v__1255_out0;
wire  [2:0] v__1256_out0;
wire  [2:0] v__1257_out0;
wire  [2:0] v__1258_out0;
wire  [2:0] v__1308_out1;
wire  [2:0] v__1444_out0;
wire  [2:0] v__1445_out0;
wire  [2:0] v__2_out0;
wire  [2:0] v__4831_out0;
wire  [2:0] v__4832_out0;
wire  [2:0] v__6536_out0;
wire  [2:0] v__841_out0;
wire  [31:0] v_32BITPRODUCT_44_out0;
wire  [31:0] v_32BITPRODUCT_6034_out0;
wire  [31:0] v_32BIT_MULTI_580_out0;
wire  [31:0] v_FLOATING_MULTI_3782_out0;
wire  [31:0] v__106_out0;
wire  [3:0] v_8BITCOUNTER_5462_out0;
wire  [3:0] v_8BITCOUNTER_6549_out0;
wire  [3:0] v_8BITCOUNTER_6550_out0;
wire  [3:0] v_BIN_2868_out0;
wire  [3:0] v_B_136_out0;
wire  [3:0] v_B_5311_out0;
wire  [3:0] v_B_567_out0;
wire  [3:0] v_C1_3397_out0;
wire  [3:0] v_C1_5082_out0;
wire  [3:0] v_C1_980_out0;
wire  [3:0] v_MUX1_1174_out0;
wire  [3:0] v_NOTUSED1_928_out0;
wire  [3:0] v_NOTUSED_4829_out0;
wire  [3:0] v_NOTUSED_5186_out0;
wire  [3:0] v_NOTUSED_6540_out0;
wire  [3:0] v_NOTUSE_1170_out0;
wire  [3:0] v_N_3755_out0;
wire  [3:0] v_RAM_ADD_BYTE0_6592_out0;
wire  [3:0] v_SEL1_2842_out0;
wire  [3:0] v_UNUSED_6616_out0;
wire  [3:0] v__1045_out0;
wire  [3:0] v__112_out1;
wire  [3:0] v__1143_out0;
wire  [3:0] v__1144_out0;
wire  [3:0] v__1175_out1;
wire  [3:0] v__1186_out0;
wire  [3:0] v__1353_out0;
wire  [3:0] v__1354_out0;
wire  [3:0] v__1448_out0;
wire  [3:0] v__1479_out1;
wire  [3:0] v__1922_out0;
wire  [3:0] v__2193_out0;
wire  [3:0] v__219_out0;
wire  [3:0] v__220_out0;
wire  [3:0] v__2213_out0;
wire  [3:0] v__2237_out0;
wire  [3:0] v__2296_out0;
wire  [3:0] v__2865_out1;
wire  [3:0] v__3452_out0;
wire  [3:0] v__3453_out0;
wire  [3:0] v__3454_out0;
wire  [3:0] v__3455_out0;
wire  [3:0] v__3456_out0;
wire  [3:0] v__3457_out0;
wire  [3:0] v__3458_out0;
wire  [3:0] v__3459_out0;
wire  [3:0] v__3460_out0;
wire  [3:0] v__3461_out0;
wire  [3:0] v__3462_out0;
wire  [3:0] v__3463_out0;
wire  [3:0] v__3464_out0;
wire  [3:0] v__3465_out0;
wire  [3:0] v__3466_out0;
wire  [3:0] v__3490_out1;
wire  [3:0] v__4276_out0;
wire  [3:0] v__4277_out0;
wire  [3:0] v__5109_out0;
wire  [3:0] v__5110_out0;
wire  [3:0] v__559_out1;
wire  [3:0] v__59_out0;
wire  [3:0] v__60_out0;
wire  [3:0] v__6554_out0;
wire  [3:0] v__6562_out0;
wire  [3:0] v__6562_out1;
wire  [4:0] v_0B00001_5193_out0;
wire  [4:0] v_A7_1328_out0;
wire  [4:0] v_B_1924_out0;
wire  [4:0] v_C10_5536_out0;
wire  [4:0] v_C14_5312_out0;
wire  [4:0] v_C1_5084_out0;
wire  [4:0] v_C1_5085_out0;
wire  [4:0] v_C4_1264_out0;
wire  [4:0] v_C8_1346_out0;
wire  [4:0] v_EXP_1188_out0;
wire  [4:0] v_EXP_1416_out0;
wire  [4:0] v_EXP_ANS_5163_out0;
wire  [4:0] v_EXP_ANS_5342_out0;
wire  [4:0] v_EXP_ANS_5443_out0;
wire  [4:0] v_EXP_ANS_6772_out0;
wire  [4:0] v_EXP_ANS_981_out0;
wire  [4:0] v_EXP_PRE_ANS_5299_out0;
wire  [4:0] v_EXP_RD_2869_out0;
wire  [4:0] v_EXP_RM_2315_out0;
wire  [4:0] v_K_1285_out0;
wire  [4:0] v_K_2838_out0;
wire  [4:0] v_MUX11_46_out0;
wire  [4:0] v_MUX12_6789_out0;
wire  [4:0] v_MUX13_6724_out0;
wire  [4:0] v_MUX4_137_out0;
wire  [4:0] v_MUX7_2189_out0;
wire  [4:0] v_OP2_EXP_1242_out0;
wire  [4:0] v_OP2_EXP_263_out0;
wire  [4:0] v_OP2_EXP_5114_out0;
wire  [4:0] v_RD_EXP_1268_out0;
wire  [4:0] v_RD_EXP_1927_out0;
wire  [4:0] v_RD_EXP_4352_out0;
wire  [4:0] v_SEL1_1421_out0;
wire  [4:0] v_SEL2_6566_out0;
wire  [4:0] v_SEL3_190_out0;
wire  [4:0] v_SEL4_2837_out0;
wire  [4:0] v_SHIFT_AMOUNT_113_out0;
wire  [4:0] v_SHIFT_AMOUNT_2302_out0;
wire  [4:0] v__1166_out0;
wire  [4:0] v__1390_out0;
wire  [4:0] v__1583_out0;
wire  [4:0] v__1584_out0;
wire  [4:0] v__2866_out0;
wire  [4:0] v__6662_out0;
wire  [4:0] v__6663_out0;
wire  [4:0] v__6664_out0;
wire  [4:0] v__6665_out0;
wire  [4:0] v__6666_out0;
wire  [4:0] v__6667_out0;
wire  [4:0] v__6668_out0;
wire  [4:0] v__6669_out0;
wire  [4:0] v__6670_out0;
wire  [4:0] v__6671_out0;
wire  [4:0] v__6672_out0;
wire  [4:0] v__6673_out0;
wire  [4:0] v__6674_out0;
wire  [4:0] v__6675_out0;
wire  [4:0] v__6676_out0;
wire  [5:0] v_A4_6704_out0;
wire  [5:0] v_A5_1286_out0;
wire  [5:0] v_A6_1931_out0;
wire  [5:0] v_C11_6781_out0;
wire  [5:0] v_C12_1029_out0;
wire  [5:0] v_C13_196_out0;
wire  [5:0] v_C9_5492_out0;
wire  [5:0] v_EXP_SUM_2864_out0;
wire  [5:0] v_MUX10_5120_out0;
wire  [5:0] v_MUX8_2238_out0;
wire  [5:0] v_MUX9_6643_out0;
wire  [5:0] v_NEG1_3398_out0;
wire  [5:0] v_NOTUSED_1317_out0;
wire  [5:0] v_XOR3_1241_out0;
wire  [5:0] v_XOR4_3417_out0;
wire  [5:0] v__1272_out0;
wire  [5:0] v__1610_out0;
wire  [5:0] v__1611_out0;
wire  [5:0] v__1612_out0;
wire  [5:0] v__1613_out0;
wire  [5:0] v__1614_out0;
wire  [5:0] v__1615_out0;
wire  [5:0] v__1616_out0;
wire  [5:0] v__1617_out0;
wire  [5:0] v__1618_out0;
wire  [5:0] v__1619_out0;
wire  [5:0] v__1620_out0;
wire  [5:0] v__1621_out0;
wire  [5:0] v__1622_out0;
wire  [5:0] v__1623_out0;
wire  [5:0] v__1624_out0;
wire  [5:0] v__1899_out1;
wire  [5:0] v__30_out0;
wire  [5:0] v__5061_out0;
wire  [5:0] v__5078_out0;
wire  [5:0] v__5079_out0;
wire  [5:0] v__50_out0;
wire  [5:0] v__5164_out0;
wire  [5:0] v__5341_out0;
wire  [6:0] v__1443_out1;
wire  [6:0] v__2296_out1;
wire  [6:0] v__330_out0;
wire  [6:0] v__3467_out0;
wire  [6:0] v__3507_out0;
wire  [6:0] v__3508_out0;
wire  [6:0] v__3509_out0;
wire  [6:0] v__3510_out0;
wire  [6:0] v__3511_out0;
wire  [6:0] v__3512_out0;
wire  [6:0] v__3513_out0;
wire  [6:0] v__3514_out0;
wire  [6:0] v__3515_out0;
wire  [6:0] v__3516_out0;
wire  [6:0] v__3517_out0;
wire  [6:0] v__3518_out0;
wire  [6:0] v__3519_out0;
wire  [6:0] v__3520_out0;
wire  [6:0] v__3521_out0;
wire  [6:0] v__37_out0;
wire  [6:0] v__62_out0;
wire  [6:0] v__63_out0;
wire  [7:0] v_C1_5063_out0;
wire  [7:0] v_C1_6547_out0;
wire  [7:0] v_C1_6623_out0;
wire  [7:0] v_MUX2_1162_out0;
wire  [7:0] v_NOTUSED2_23_out0;
wire  [7:0] v_NOTUSED_331_out0;
wire  [7:0] v_NOTUSED_35_out0;
wire  [7:0] v_NOTUSED_5198_out0;
wire  [7:0] v_OUT_1480_out0;
wire  [7:0] v_RECEIVERSTREAM_3751_out0;
wire  [7:0] v_RECEIVER_STREAM_276_out0;
wire  [7:0] v_RECEIVER_STREAM_6544_out0;
wire  [7:0] v_RECEIVER_stream_5189_out0;
wire  [7:0] v_REGISTER_TRANSMIT_DATA_6031_out0;
wire  [7:0] v_TRANSMISSION_DATA_1327_out0;
wire  [7:0] v_TRANSMIT_DATA_39_out0;
wire  [7:0] v__1186_out1;
wire  [7:0] v__1259_out0;
wire  [7:0] v__1259_out1;
wire  [7:0] v__1308_out0;
wire  [7:0] v__1310_out0;
wire  [7:0] v__1311_out0;
wire  [7:0] v__1482_out0;
wire  [7:0] v__1524_out0;
wire  [7:0] v__1524_out1;
wire  [7:0] v__2176_out0;
wire  [7:0] v__2177_out0;
wire  [7:0] v__2318_out0;
wire  [7:0] v__2319_out0;
wire  [7:0] v__2320_out0;
wire  [7:0] v__2321_out0;
wire  [7:0] v__2322_out0;
wire  [7:0] v__2323_out0;
wire  [7:0] v__2324_out0;
wire  [7:0] v__2325_out0;
wire  [7:0] v__2326_out0;
wire  [7:0] v__2327_out0;
wire  [7:0] v__2328_out0;
wire  [7:0] v__2329_out0;
wire  [7:0] v__2330_out0;
wire  [7:0] v__2331_out0;
wire  [7:0] v__2332_out0;
wire  [7:0] v__308_out0;
wire  [7:0] v__4270_out0;
wire  [7:0] v__4270_out1;
wire  [7:0] v__4274_out0;
wire  [7:0] v__5347_out0;
wire  [7:0] v__5480_out0;
wire  [7:0] v__5480_out1;
wire  [7:0] v__6793_out0;
wire  [7:0] v__6794_out0;
wire  [7:0] v_split_214_out0;
wire  [7:0] v_split_214_out1;
wire  [8:0] v_SEL6_1948_out0;
wire  [8:0] v__1386_out0;
wire  [8:0] v__2211_out0;
wire  [8:0] v__227_out0;
wire  [8:0] v__228_out0;
wire  [8:0] v__24_out0;
wire  [8:0] v__3400_out0;
wire  [8:0] v__3401_out0;
wire  [8:0] v__3402_out0;
wire  [8:0] v__3403_out0;
wire  [8:0] v__3404_out0;
wire  [8:0] v__3405_out0;
wire  [8:0] v__3406_out0;
wire  [8:0] v__3407_out0;
wire  [8:0] v__3408_out0;
wire  [8:0] v__3409_out0;
wire  [8:0] v__3410_out0;
wire  [8:0] v__3411_out0;
wire  [8:0] v__3412_out0;
wire  [8:0] v__3413_out0;
wire  [8:0] v__3414_out0;
wire  [8:0] v__3785_out0;
wire  [8:0] v__6678_out1;
wire  [9:0] v_MUX4_5103_out0;
wire  [9:0] v_MUX6_5100_out0;
wire  [9:0] v_OP2_SIG_6556_out0;
wire  [9:0] v_RD_SIG_865_out0;
wire  [9:0] v_SEL4_5525_out0;
wire  [9:0] v_SEL5_4314_out0;
wire  [9:0] v_SEL6_53_out0;
wire  [9:0] v_SEL9_6774_out0;
wire  [9:0] v_SIG_ANS_1139_out0;
wire  [9:0] v_SIG_ANS_1593_out0;
wire  [9:0] v_SIG_ANS_213_out0;
wire  [9:0] v_SIG_ANS_5077_out0;
wire  [9:0] v_SIG_RD_5561_out0;
wire  [9:0] v_SIG_RM_864_out0;
wire  [9:0] v__1291_out0;
wire  [9:0] v__1899_out0;
wire  [9:0] v__1905_out1;
wire  [9:0] v__206_out0;
wire  [9:0] v__207_out0;
wire  [9:0] v__2844_out0;
wire  [9:0] v__2845_out0;
wire  [9:0] v__2846_out0;
wire  [9:0] v__2847_out0;
wire  [9:0] v__2848_out0;
wire  [9:0] v__2849_out0;
wire  [9:0] v__2850_out0;
wire  [9:0] v__2851_out0;
wire  [9:0] v__2852_out0;
wire  [9:0] v__2853_out0;
wire  [9:0] v__2854_out0;
wire  [9:0] v__2855_out0;
wire  [9:0] v__2856_out0;
wire  [9:0] v__2857_out0;
wire  [9:0] v__2858_out0;
wire  [9:0] v__4272_out0;
wire  [9:0] v__5303_out0;
wire  [9:0] v__5316_out0;
wire v_0_1475_out0;
wire v_0_5269_out0;
wire v_1_1860_out0;
wire v_2_3472_out0;
wire v_2_862_out0;
wire v_3_6711_out0;
wire v_9_203_out0;
wire v_9_6712_out0;
wire v_9_6713_out0;
wire v_9_834_out0;
wire v_9_835_out0;
wire v_A1_1547_out1;
wire v_A1_1879_out1;
wire v_A1_3446_out1;
wire v_A1_5433_out1;
wire v_A4_5526_out1;
wire v_A4_6704_out1;
wire v_A5_1286_out1;
wire v_A5_929_out1;
wire v_A6_1931_out1;
wire v_A6_5152_out1;
wire v_A7_1328_out1;
wire v_A8_5490_out1;
wire v_ADC_5119_out0;
wire v_ADC_6710_out0;
wire v_ADC_889_out0;
wire v_ADD_2179_out0;
wire v_ADD_5509_out0;
wire v_AND_1880_out0;
wire v_AND_6681_out0;
wire v_ASR_4308_out0;
wire v_ASR_5107_out0;
wire v_ASR_5199_out0;
wire v_ASR_6755_out0;
wire v_BIT10_3441_out0;
wire v_BIT_1135_out0;
wire v_BIT_3396_out0;
wire v_BIT_STREAM_IN_7_out0;
wire v_BYTE1_comp1_1189_out0;
wire v_BYTE2_COMP8_3781_out0;
wire v_BYTERECEIVED_5511_out0;
wire v_BYTE_READY_1393_out0;
wire v_BYTE_READY_2239_out0;
wire v_BYTE_READY_3447_out0;
wire v_BYTE_READY_5195_out0;
wire v_BYTE_READY_5498_out0;
wire v_BYTE_READY_RX_4826_out0;
wire v_C10_888_out0;
wire v_C12_565_out0;
wire v_C14_822_out0;
wire v_C1_211_out0;
wire v_C1_293_out0;
wire v_C1_4338_out0;
wire v_C1_5058_out0;
wire v_C1_5309_out0;
wire v_C3_2314_out0;
wire v_C4_5227_out0;
wire v_C5_6541_out0;
wire v_C6_5086_out0;
wire v_C7_1108_out0;
wire v_C9_1477_out0;
wire v_CARRY_2373_out0;
wire v_CARRY_2374_out0;
wire v_CARRY_2375_out0;
wire v_CARRY_2376_out0;
wire v_CARRY_2377_out0;
wire v_CARRY_2378_out0;
wire v_CARRY_2379_out0;
wire v_CARRY_2380_out0;
wire v_CARRY_2381_out0;
wire v_CARRY_2382_out0;
wire v_CARRY_2383_out0;
wire v_CARRY_2384_out0;
wire v_CARRY_2385_out0;
wire v_CARRY_2386_out0;
wire v_CARRY_2387_out0;
wire v_CARRY_2388_out0;
wire v_CARRY_2389_out0;
wire v_CARRY_2390_out0;
wire v_CARRY_2391_out0;
wire v_CARRY_2392_out0;
wire v_CARRY_2393_out0;
wire v_CARRY_2394_out0;
wire v_CARRY_2395_out0;
wire v_CARRY_2396_out0;
wire v_CARRY_2397_out0;
wire v_CARRY_2398_out0;
wire v_CARRY_2399_out0;
wire v_CARRY_2400_out0;
wire v_CARRY_2401_out0;
wire v_CARRY_2402_out0;
wire v_CARRY_2403_out0;
wire v_CARRY_2404_out0;
wire v_CARRY_2405_out0;
wire v_CARRY_2406_out0;
wire v_CARRY_2407_out0;
wire v_CARRY_2408_out0;
wire v_CARRY_2409_out0;
wire v_CARRY_2410_out0;
wire v_CARRY_2411_out0;
wire v_CARRY_2412_out0;
wire v_CARRY_2413_out0;
wire v_CARRY_2414_out0;
wire v_CARRY_2415_out0;
wire v_CARRY_2416_out0;
wire v_CARRY_2417_out0;
wire v_CARRY_2418_out0;
wire v_CARRY_2419_out0;
wire v_CARRY_2420_out0;
wire v_CARRY_2421_out0;
wire v_CARRY_2422_out0;
wire v_CARRY_2423_out0;
wire v_CARRY_2424_out0;
wire v_CARRY_2425_out0;
wire v_CARRY_2426_out0;
wire v_CARRY_2427_out0;
wire v_CARRY_2428_out0;
wire v_CARRY_2429_out0;
wire v_CARRY_2430_out0;
wire v_CARRY_2431_out0;
wire v_CARRY_2432_out0;
wire v_CARRY_2433_out0;
wire v_CARRY_2434_out0;
wire v_CARRY_2435_out0;
wire v_CARRY_2436_out0;
wire v_CARRY_2437_out0;
wire v_CARRY_2438_out0;
wire v_CARRY_2439_out0;
wire v_CARRY_2440_out0;
wire v_CARRY_2441_out0;
wire v_CARRY_2442_out0;
wire v_CARRY_2443_out0;
wire v_CARRY_2444_out0;
wire v_CARRY_2445_out0;
wire v_CARRY_2446_out0;
wire v_CARRY_2447_out0;
wire v_CARRY_2448_out0;
wire v_CARRY_2449_out0;
wire v_CARRY_2450_out0;
wire v_CARRY_2451_out0;
wire v_CARRY_2452_out0;
wire v_CARRY_2453_out0;
wire v_CARRY_2454_out0;
wire v_CARRY_2455_out0;
wire v_CARRY_2456_out0;
wire v_CARRY_2457_out0;
wire v_CARRY_2458_out0;
wire v_CARRY_2459_out0;
wire v_CARRY_2460_out0;
wire v_CARRY_2461_out0;
wire v_CARRY_2462_out0;
wire v_CARRY_2463_out0;
wire v_CARRY_2464_out0;
wire v_CARRY_2465_out0;
wire v_CARRY_2466_out0;
wire v_CARRY_2467_out0;
wire v_CARRY_2468_out0;
wire v_CARRY_2469_out0;
wire v_CARRY_2470_out0;
wire v_CARRY_2471_out0;
wire v_CARRY_2472_out0;
wire v_CARRY_2473_out0;
wire v_CARRY_2474_out0;
wire v_CARRY_2475_out0;
wire v_CARRY_2476_out0;
wire v_CARRY_2477_out0;
wire v_CARRY_2478_out0;
wire v_CARRY_2479_out0;
wire v_CARRY_2480_out0;
wire v_CARRY_2481_out0;
wire v_CARRY_2482_out0;
wire v_CARRY_2483_out0;
wire v_CARRY_2484_out0;
wire v_CARRY_2485_out0;
wire v_CARRY_2486_out0;
wire v_CARRY_2487_out0;
wire v_CARRY_2488_out0;
wire v_CARRY_2489_out0;
wire v_CARRY_2490_out0;
wire v_CARRY_2491_out0;
wire v_CARRY_2492_out0;
wire v_CARRY_2493_out0;
wire v_CARRY_2494_out0;
wire v_CARRY_2495_out0;
wire v_CARRY_2496_out0;
wire v_CARRY_2497_out0;
wire v_CARRY_2498_out0;
wire v_CARRY_2499_out0;
wire v_CARRY_2500_out0;
wire v_CARRY_2501_out0;
wire v_CARRY_2502_out0;
wire v_CARRY_2503_out0;
wire v_CARRY_2504_out0;
wire v_CARRY_2505_out0;
wire v_CARRY_2506_out0;
wire v_CARRY_2507_out0;
wire v_CARRY_2508_out0;
wire v_CARRY_2509_out0;
wire v_CARRY_2510_out0;
wire v_CARRY_2511_out0;
wire v_CARRY_2512_out0;
wire v_CARRY_2513_out0;
wire v_CARRY_2514_out0;
wire v_CARRY_2515_out0;
wire v_CARRY_2516_out0;
wire v_CARRY_2517_out0;
wire v_CARRY_2518_out0;
wire v_CARRY_2519_out0;
wire v_CARRY_2520_out0;
wire v_CARRY_2521_out0;
wire v_CARRY_2522_out0;
wire v_CARRY_2523_out0;
wire v_CARRY_2524_out0;
wire v_CARRY_2525_out0;
wire v_CARRY_2526_out0;
wire v_CARRY_2527_out0;
wire v_CARRY_2528_out0;
wire v_CARRY_2529_out0;
wire v_CARRY_2530_out0;
wire v_CARRY_2531_out0;
wire v_CARRY_2532_out0;
wire v_CARRY_2533_out0;
wire v_CARRY_2534_out0;
wire v_CARRY_2535_out0;
wire v_CARRY_2536_out0;
wire v_CARRY_2537_out0;
wire v_CARRY_2538_out0;
wire v_CARRY_2539_out0;
wire v_CARRY_2540_out0;
wire v_CARRY_2541_out0;
wire v_CARRY_2542_out0;
wire v_CARRY_2543_out0;
wire v_CARRY_2544_out0;
wire v_CARRY_2545_out0;
wire v_CARRY_2546_out0;
wire v_CARRY_2547_out0;
wire v_CARRY_2548_out0;
wire v_CARRY_2549_out0;
wire v_CARRY_2550_out0;
wire v_CARRY_2551_out0;
wire v_CARRY_2552_out0;
wire v_CARRY_2553_out0;
wire v_CARRY_2554_out0;
wire v_CARRY_2555_out0;
wire v_CARRY_2556_out0;
wire v_CARRY_2557_out0;
wire v_CARRY_2558_out0;
wire v_CARRY_2559_out0;
wire v_CARRY_2560_out0;
wire v_CARRY_2561_out0;
wire v_CARRY_2562_out0;
wire v_CARRY_2563_out0;
wire v_CARRY_2564_out0;
wire v_CARRY_2565_out0;
wire v_CARRY_2566_out0;
wire v_CARRY_2567_out0;
wire v_CARRY_2568_out0;
wire v_CARRY_2569_out0;
wire v_CARRY_2570_out0;
wire v_CARRY_2571_out0;
wire v_CARRY_2572_out0;
wire v_CARRY_2573_out0;
wire v_CARRY_2574_out0;
wire v_CARRY_2575_out0;
wire v_CARRY_2576_out0;
wire v_CARRY_2577_out0;
wire v_CARRY_2578_out0;
wire v_CARRY_2579_out0;
wire v_CARRY_2580_out0;
wire v_CARRY_2581_out0;
wire v_CARRY_2582_out0;
wire v_CARRY_2583_out0;
wire v_CARRY_2584_out0;
wire v_CARRY_2585_out0;
wire v_CARRY_2586_out0;
wire v_CARRY_2587_out0;
wire v_CARRY_2588_out0;
wire v_CARRY_2589_out0;
wire v_CARRY_2590_out0;
wire v_CARRY_2591_out0;
wire v_CARRY_2592_out0;
wire v_CARRY_2593_out0;
wire v_CARRY_2594_out0;
wire v_CARRY_2595_out0;
wire v_CARRY_2596_out0;
wire v_CARRY_2597_out0;
wire v_CARRY_2598_out0;
wire v_CARRY_2599_out0;
wire v_CARRY_2600_out0;
wire v_CARRY_2601_out0;
wire v_CARRY_2602_out0;
wire v_CARRY_2603_out0;
wire v_CARRY_2604_out0;
wire v_CARRY_2605_out0;
wire v_CARRY_2606_out0;
wire v_CARRY_2607_out0;
wire v_CARRY_2608_out0;
wire v_CARRY_2609_out0;
wire v_CARRY_2610_out0;
wire v_CARRY_2611_out0;
wire v_CARRY_2612_out0;
wire v_CARRY_2613_out0;
wire v_CARRY_2614_out0;
wire v_CARRY_2615_out0;
wire v_CARRY_2616_out0;
wire v_CARRY_2617_out0;
wire v_CARRY_2618_out0;
wire v_CARRY_2619_out0;
wire v_CARRY_2620_out0;
wire v_CARRY_2621_out0;
wire v_CARRY_2622_out0;
wire v_CARRY_2623_out0;
wire v_CARRY_2624_out0;
wire v_CARRY_2625_out0;
wire v_CARRY_2626_out0;
wire v_CARRY_2627_out0;
wire v_CARRY_2628_out0;
wire v_CARRY_2629_out0;
wire v_CARRY_2630_out0;
wire v_CARRY_2631_out0;
wire v_CARRY_2632_out0;
wire v_CARRY_2633_out0;
wire v_CARRY_2634_out0;
wire v_CARRY_2635_out0;
wire v_CARRY_2636_out0;
wire v_CARRY_2637_out0;
wire v_CARRY_2638_out0;
wire v_CARRY_2639_out0;
wire v_CARRY_2640_out0;
wire v_CARRY_2641_out0;
wire v_CARRY_2642_out0;
wire v_CARRY_2643_out0;
wire v_CARRY_2644_out0;
wire v_CARRY_2645_out0;
wire v_CARRY_2646_out0;
wire v_CARRY_2647_out0;
wire v_CARRY_2648_out0;
wire v_CARRY_2649_out0;
wire v_CARRY_2650_out0;
wire v_CARRY_2651_out0;
wire v_CARRY_2652_out0;
wire v_CARRY_2653_out0;
wire v_CARRY_2654_out0;
wire v_CARRY_2655_out0;
wire v_CARRY_2656_out0;
wire v_CARRY_2657_out0;
wire v_CARRY_2658_out0;
wire v_CARRY_2659_out0;
wire v_CARRY_2660_out0;
wire v_CARRY_2661_out0;
wire v_CARRY_2662_out0;
wire v_CARRY_2663_out0;
wire v_CARRY_2664_out0;
wire v_CARRY_2665_out0;
wire v_CARRY_2666_out0;
wire v_CARRY_2667_out0;
wire v_CARRY_2668_out0;
wire v_CARRY_2669_out0;
wire v_CARRY_2670_out0;
wire v_CARRY_2671_out0;
wire v_CARRY_2672_out0;
wire v_CARRY_2673_out0;
wire v_CARRY_2674_out0;
wire v_CARRY_2675_out0;
wire v_CARRY_2676_out0;
wire v_CARRY_2677_out0;
wire v_CARRY_2678_out0;
wire v_CARRY_2679_out0;
wire v_CARRY_2680_out0;
wire v_CARRY_2681_out0;
wire v_CARRY_2682_out0;
wire v_CARRY_2683_out0;
wire v_CARRY_2684_out0;
wire v_CARRY_2685_out0;
wire v_CARRY_2686_out0;
wire v_CARRY_2687_out0;
wire v_CARRY_2688_out0;
wire v_CARRY_2689_out0;
wire v_CARRY_2690_out0;
wire v_CARRY_2691_out0;
wire v_CARRY_2692_out0;
wire v_CARRY_2693_out0;
wire v_CARRY_2694_out0;
wire v_CARRY_2695_out0;
wire v_CARRY_2696_out0;
wire v_CARRY_2697_out0;
wire v_CARRY_2698_out0;
wire v_CARRY_2699_out0;
wire v_CARRY_2700_out0;
wire v_CARRY_2701_out0;
wire v_CARRY_2702_out0;
wire v_CARRY_2703_out0;
wire v_CARRY_2704_out0;
wire v_CARRY_2705_out0;
wire v_CARRY_2706_out0;
wire v_CARRY_2707_out0;
wire v_CARRY_2708_out0;
wire v_CARRY_2709_out0;
wire v_CARRY_2710_out0;
wire v_CARRY_2711_out0;
wire v_CARRY_2712_out0;
wire v_CARRY_2713_out0;
wire v_CARRY_2714_out0;
wire v_CARRY_2715_out0;
wire v_CARRY_2716_out0;
wire v_CARRY_2717_out0;
wire v_CARRY_2718_out0;
wire v_CARRY_2719_out0;
wire v_CARRY_2720_out0;
wire v_CARRY_2721_out0;
wire v_CARRY_2722_out0;
wire v_CARRY_2723_out0;
wire v_CARRY_2724_out0;
wire v_CARRY_2725_out0;
wire v_CARRY_2726_out0;
wire v_CARRY_2727_out0;
wire v_CARRY_2728_out0;
wire v_CARRY_2729_out0;
wire v_CARRY_2730_out0;
wire v_CARRY_2731_out0;
wire v_CARRY_2732_out0;
wire v_CARRY_2733_out0;
wire v_CARRY_2734_out0;
wire v_CARRY_2735_out0;
wire v_CARRY_2736_out0;
wire v_CARRY_2737_out0;
wire v_CARRY_2738_out0;
wire v_CARRY_2739_out0;
wire v_CARRY_2740_out0;
wire v_CARRY_2741_out0;
wire v_CARRY_2742_out0;
wire v_CARRY_2743_out0;
wire v_CARRY_2744_out0;
wire v_CARRY_2745_out0;
wire v_CARRY_2746_out0;
wire v_CARRY_2747_out0;
wire v_CARRY_2748_out0;
wire v_CARRY_2749_out0;
wire v_CARRY_2750_out0;
wire v_CARRY_2751_out0;
wire v_CARRY_2752_out0;
wire v_CARRY_2753_out0;
wire v_CARRY_2754_out0;
wire v_CARRY_2755_out0;
wire v_CARRY_2756_out0;
wire v_CARRY_2757_out0;
wire v_CARRY_2758_out0;
wire v_CARRY_2759_out0;
wire v_CARRY_2760_out0;
wire v_CARRY_2761_out0;
wire v_CARRY_2762_out0;
wire v_CARRY_2763_out0;
wire v_CARRY_2764_out0;
wire v_CARRY_2765_out0;
wire v_CARRY_2766_out0;
wire v_CARRY_2767_out0;
wire v_CARRY_2768_out0;
wire v_CARRY_2769_out0;
wire v_CARRY_2770_out0;
wire v_CARRY_2771_out0;
wire v_CARRY_2772_out0;
wire v_CARRY_2773_out0;
wire v_CARRY_2774_out0;
wire v_CARRY_2775_out0;
wire v_CARRY_2776_out0;
wire v_CARRY_2777_out0;
wire v_CARRY_2778_out0;
wire v_CARRY_2779_out0;
wire v_CARRY_2780_out0;
wire v_CARRY_2781_out0;
wire v_CARRY_2782_out0;
wire v_CARRY_2783_out0;
wire v_CARRY_2784_out0;
wire v_CARRY_2785_out0;
wire v_CARRY_2786_out0;
wire v_CARRY_2787_out0;
wire v_CARRY_2788_out0;
wire v_CARRY_2789_out0;
wire v_CARRY_2790_out0;
wire v_CARRY_2791_out0;
wire v_CARRY_2792_out0;
wire v_CARRY_2793_out0;
wire v_CARRY_2794_out0;
wire v_CARRY_2795_out0;
wire v_CARRY_2796_out0;
wire v_CARRY_2797_out0;
wire v_CARRY_2798_out0;
wire v_CARRY_2799_out0;
wire v_CARRY_2800_out0;
wire v_CARRY_2801_out0;
wire v_CARRY_2802_out0;
wire v_CARRY_2803_out0;
wire v_CARRY_2804_out0;
wire v_CARRY_2805_out0;
wire v_CARRY_2806_out0;
wire v_CARRY_2807_out0;
wire v_CARRY_2808_out0;
wire v_CARRY_2809_out0;
wire v_CARRY_2810_out0;
wire v_CARRY_2811_out0;
wire v_CARRY_2812_out0;
wire v_CARRY_2813_out0;
wire v_CARRY_2814_out0;
wire v_CARRY_2815_out0;
wire v_CARRY_2816_out0;
wire v_CARRY_2817_out0;
wire v_CARRY_2818_out0;
wire v_CARRY_2819_out0;
wire v_CARRY_2820_out0;
wire v_CARRY_2821_out0;
wire v_CARRY_2822_out0;
wire v_CARRY_2823_out0;
wire v_CARRY_2824_out0;
wire v_CARRY_2825_out0;
wire v_CARRY_2826_out0;
wire v_CARRY_2827_out0;
wire v_CARRY_2828_out0;
wire v_CARRY_2829_out0;
wire v_CARRY_2830_out0;
wire v_CARRY_2831_out0;
wire v_CARRY_2832_out0;
wire v_CARRY_2833_out0;
wire v_CARRY_2834_out0;
wire v_CARRY_2835_out0;
wire v_CARRY_2836_out0;
wire v_CIN_4833_out0;
wire v_CIN_4834_out0;
wire v_CIN_4835_out0;
wire v_CIN_4836_out0;
wire v_CIN_4837_out0;
wire v_CIN_4838_out0;
wire v_CIN_4839_out0;
wire v_CIN_4840_out0;
wire v_CIN_4841_out0;
wire v_CIN_4842_out0;
wire v_CIN_4843_out0;
wire v_CIN_4844_out0;
wire v_CIN_4845_out0;
wire v_CIN_4846_out0;
wire v_CIN_4847_out0;
wire v_CIN_4848_out0;
wire v_CIN_4849_out0;
wire v_CIN_4850_out0;
wire v_CIN_4851_out0;
wire v_CIN_4852_out0;
wire v_CIN_4853_out0;
wire v_CIN_4854_out0;
wire v_CIN_4855_out0;
wire v_CIN_4856_out0;
wire v_CIN_4857_out0;
wire v_CIN_4858_out0;
wire v_CIN_4859_out0;
wire v_CIN_4860_out0;
wire v_CIN_4861_out0;
wire v_CIN_4862_out0;
wire v_CIN_4863_out0;
wire v_CIN_4864_out0;
wire v_CIN_4865_out0;
wire v_CIN_4866_out0;
wire v_CIN_4867_out0;
wire v_CIN_4868_out0;
wire v_CIN_4869_out0;
wire v_CIN_4870_out0;
wire v_CIN_4871_out0;
wire v_CIN_4872_out0;
wire v_CIN_4873_out0;
wire v_CIN_4874_out0;
wire v_CIN_4875_out0;
wire v_CIN_4876_out0;
wire v_CIN_4877_out0;
wire v_CIN_4878_out0;
wire v_CIN_4879_out0;
wire v_CIN_4880_out0;
wire v_CIN_4881_out0;
wire v_CIN_4882_out0;
wire v_CIN_4883_out0;
wire v_CIN_4884_out0;
wire v_CIN_4885_out0;
wire v_CIN_4886_out0;
wire v_CIN_4887_out0;
wire v_CIN_4888_out0;
wire v_CIN_4889_out0;
wire v_CIN_4890_out0;
wire v_CIN_4891_out0;
wire v_CIN_4892_out0;
wire v_CIN_4893_out0;
wire v_CIN_4894_out0;
wire v_CIN_4895_out0;
wire v_CIN_4896_out0;
wire v_CIN_4897_out0;
wire v_CIN_4898_out0;
wire v_CIN_4899_out0;
wire v_CIN_4900_out0;
wire v_CIN_4901_out0;
wire v_CIN_4902_out0;
wire v_CIN_4903_out0;
wire v_CIN_4904_out0;
wire v_CIN_4905_out0;
wire v_CIN_4906_out0;
wire v_CIN_4907_out0;
wire v_CIN_4908_out0;
wire v_CIN_4909_out0;
wire v_CIN_4910_out0;
wire v_CIN_4911_out0;
wire v_CIN_4912_out0;
wire v_CIN_4913_out0;
wire v_CIN_4914_out0;
wire v_CIN_4915_out0;
wire v_CIN_4916_out0;
wire v_CIN_4917_out0;
wire v_CIN_4918_out0;
wire v_CIN_4919_out0;
wire v_CIN_4920_out0;
wire v_CIN_4921_out0;
wire v_CIN_4922_out0;
wire v_CIN_4923_out0;
wire v_CIN_4924_out0;
wire v_CIN_4925_out0;
wire v_CIN_4926_out0;
wire v_CIN_4927_out0;
wire v_CIN_4928_out0;
wire v_CIN_4929_out0;
wire v_CIN_4930_out0;
wire v_CIN_4931_out0;
wire v_CIN_4932_out0;
wire v_CIN_4933_out0;
wire v_CIN_4934_out0;
wire v_CIN_4935_out0;
wire v_CIN_4936_out0;
wire v_CIN_4937_out0;
wire v_CIN_4938_out0;
wire v_CIN_4939_out0;
wire v_CIN_4940_out0;
wire v_CIN_4941_out0;
wire v_CIN_4942_out0;
wire v_CIN_4943_out0;
wire v_CIN_4944_out0;
wire v_CIN_4945_out0;
wire v_CIN_4946_out0;
wire v_CIN_4947_out0;
wire v_CIN_4948_out0;
wire v_CIN_4949_out0;
wire v_CIN_4950_out0;
wire v_CIN_4951_out0;
wire v_CIN_4952_out0;
wire v_CIN_4953_out0;
wire v_CIN_4954_out0;
wire v_CIN_4955_out0;
wire v_CIN_4956_out0;
wire v_CIN_4957_out0;
wire v_CIN_4958_out0;
wire v_CIN_4959_out0;
wire v_CIN_4960_out0;
wire v_CIN_4961_out0;
wire v_CIN_4962_out0;
wire v_CIN_4963_out0;
wire v_CIN_4964_out0;
wire v_CIN_4965_out0;
wire v_CIN_4966_out0;
wire v_CIN_4967_out0;
wire v_CIN_4968_out0;
wire v_CIN_4969_out0;
wire v_CIN_4970_out0;
wire v_CIN_4971_out0;
wire v_CIN_4972_out0;
wire v_CIN_4973_out0;
wire v_CIN_4974_out0;
wire v_CIN_4975_out0;
wire v_CIN_4976_out0;
wire v_CIN_4977_out0;
wire v_CIN_4978_out0;
wire v_CIN_4979_out0;
wire v_CIN_4980_out0;
wire v_CIN_4981_out0;
wire v_CIN_4982_out0;
wire v_CIN_4983_out0;
wire v_CIN_4984_out0;
wire v_CIN_4985_out0;
wire v_CIN_4986_out0;
wire v_CIN_4987_out0;
wire v_CIN_4988_out0;
wire v_CIN_4989_out0;
wire v_CIN_4990_out0;
wire v_CIN_4991_out0;
wire v_CIN_4992_out0;
wire v_CIN_4993_out0;
wire v_CIN_4994_out0;
wire v_CIN_4995_out0;
wire v_CIN_4996_out0;
wire v_CIN_4997_out0;
wire v_CIN_4998_out0;
wire v_CIN_4999_out0;
wire v_CIN_5000_out0;
wire v_CIN_5001_out0;
wire v_CIN_5002_out0;
wire v_CIN_5003_out0;
wire v_CIN_5004_out0;
wire v_CIN_5005_out0;
wire v_CIN_5006_out0;
wire v_CIN_5007_out0;
wire v_CIN_5008_out0;
wire v_CIN_5009_out0;
wire v_CIN_5010_out0;
wire v_CIN_5011_out0;
wire v_CIN_5012_out0;
wire v_CIN_5013_out0;
wire v_CIN_5014_out0;
wire v_CIN_5015_out0;
wire v_CIN_5016_out0;
wire v_CIN_5017_out0;
wire v_CIN_5018_out0;
wire v_CIN_5019_out0;
wire v_CIN_5020_out0;
wire v_CIN_5021_out0;
wire v_CIN_5022_out0;
wire v_CIN_5023_out0;
wire v_CIN_5024_out0;
wire v_CIN_5025_out0;
wire v_CIN_5026_out0;
wire v_CIN_5027_out0;
wire v_CIN_5028_out0;
wire v_CIN_5029_out0;
wire v_CIN_5030_out0;
wire v_CIN_5031_out0;
wire v_CIN_5032_out0;
wire v_CIN_5033_out0;
wire v_CIN_5034_out0;
wire v_CIN_5035_out0;
wire v_CIN_5036_out0;
wire v_CIN_5037_out0;
wire v_CIN_5038_out0;
wire v_CIN_5039_out0;
wire v_CIN_5040_out0;
wire v_CIN_5041_out0;
wire v_CIN_5042_out0;
wire v_CIN_5043_out0;
wire v_CIN_5044_out0;
wire v_CIN_5045_out0;
wire v_CIN_5046_out0;
wire v_CIN_5047_out0;
wire v_CIN_5048_out0;
wire v_CIN_5049_out0;
wire v_CIN_5050_out0;
wire v_CIN_5051_out0;
wire v_CIN_5052_out0;
wire v_CIN_5053_out0;
wire v_CIN_5054_out0;
wire v_CIN_5055_out0;
wire v_CIN_5056_out0;
wire v_CMP_1855_out0;
wire v_CMP_4255_out0;
wire v_CMP_6707_out0;
wire v_COUT_1330_out0;
wire v_COUT_1898_out0;
wire v_COUT_333_out0;
wire v_COUT_334_out0;
wire v_COUT_335_out0;
wire v_COUT_336_out0;
wire v_COUT_337_out0;
wire v_COUT_338_out0;
wire v_COUT_339_out0;
wire v_COUT_340_out0;
wire v_COUT_341_out0;
wire v_COUT_342_out0;
wire v_COUT_343_out0;
wire v_COUT_344_out0;
wire v_COUT_345_out0;
wire v_COUT_346_out0;
wire v_COUT_347_out0;
wire v_COUT_348_out0;
wire v_COUT_349_out0;
wire v_COUT_350_out0;
wire v_COUT_351_out0;
wire v_COUT_352_out0;
wire v_COUT_353_out0;
wire v_COUT_354_out0;
wire v_COUT_355_out0;
wire v_COUT_356_out0;
wire v_COUT_357_out0;
wire v_COUT_358_out0;
wire v_COUT_359_out0;
wire v_COUT_360_out0;
wire v_COUT_361_out0;
wire v_COUT_362_out0;
wire v_COUT_363_out0;
wire v_COUT_364_out0;
wire v_COUT_365_out0;
wire v_COUT_366_out0;
wire v_COUT_367_out0;
wire v_COUT_368_out0;
wire v_COUT_369_out0;
wire v_COUT_36_out0;
wire v_COUT_370_out0;
wire v_COUT_371_out0;
wire v_COUT_372_out0;
wire v_COUT_373_out0;
wire v_COUT_374_out0;
wire v_COUT_375_out0;
wire v_COUT_376_out0;
wire v_COUT_377_out0;
wire v_COUT_378_out0;
wire v_COUT_379_out0;
wire v_COUT_380_out0;
wire v_COUT_381_out0;
wire v_COUT_382_out0;
wire v_COUT_383_out0;
wire v_COUT_384_out0;
wire v_COUT_385_out0;
wire v_COUT_386_out0;
wire v_COUT_387_out0;
wire v_COUT_388_out0;
wire v_COUT_389_out0;
wire v_COUT_390_out0;
wire v_COUT_391_out0;
wire v_COUT_392_out0;
wire v_COUT_393_out0;
wire v_COUT_394_out0;
wire v_COUT_395_out0;
wire v_COUT_396_out0;
wire v_COUT_397_out0;
wire v_COUT_398_out0;
wire v_COUT_399_out0;
wire v_COUT_400_out0;
wire v_COUT_401_out0;
wire v_COUT_402_out0;
wire v_COUT_403_out0;
wire v_COUT_404_out0;
wire v_COUT_405_out0;
wire v_COUT_406_out0;
wire v_COUT_407_out0;
wire v_COUT_408_out0;
wire v_COUT_409_out0;
wire v_COUT_410_out0;
wire v_COUT_411_out0;
wire v_COUT_412_out0;
wire v_COUT_413_out0;
wire v_COUT_414_out0;
wire v_COUT_415_out0;
wire v_COUT_416_out0;
wire v_COUT_417_out0;
wire v_COUT_418_out0;
wire v_COUT_419_out0;
wire v_COUT_420_out0;
wire v_COUT_421_out0;
wire v_COUT_422_out0;
wire v_COUT_423_out0;
wire v_COUT_424_out0;
wire v_COUT_425_out0;
wire v_COUT_426_out0;
wire v_COUT_427_out0;
wire v_COUT_428_out0;
wire v_COUT_429_out0;
wire v_COUT_430_out0;
wire v_COUT_431_out0;
wire v_COUT_432_out0;
wire v_COUT_433_out0;
wire v_COUT_434_out0;
wire v_COUT_435_out0;
wire v_COUT_436_out0;
wire v_COUT_437_out0;
wire v_COUT_438_out0;
wire v_COUT_439_out0;
wire v_COUT_440_out0;
wire v_COUT_441_out0;
wire v_COUT_442_out0;
wire v_COUT_443_out0;
wire v_COUT_444_out0;
wire v_COUT_445_out0;
wire v_COUT_446_out0;
wire v_COUT_447_out0;
wire v_COUT_448_out0;
wire v_COUT_449_out0;
wire v_COUT_450_out0;
wire v_COUT_451_out0;
wire v_COUT_452_out0;
wire v_COUT_453_out0;
wire v_COUT_454_out0;
wire v_COUT_455_out0;
wire v_COUT_456_out0;
wire v_COUT_457_out0;
wire v_COUT_458_out0;
wire v_COUT_459_out0;
wire v_COUT_460_out0;
wire v_COUT_461_out0;
wire v_COUT_462_out0;
wire v_COUT_463_out0;
wire v_COUT_464_out0;
wire v_COUT_465_out0;
wire v_COUT_466_out0;
wire v_COUT_467_out0;
wire v_COUT_468_out0;
wire v_COUT_469_out0;
wire v_COUT_470_out0;
wire v_COUT_471_out0;
wire v_COUT_472_out0;
wire v_COUT_473_out0;
wire v_COUT_474_out0;
wire v_COUT_475_out0;
wire v_COUT_476_out0;
wire v_COUT_477_out0;
wire v_COUT_478_out0;
wire v_COUT_479_out0;
wire v_COUT_480_out0;
wire v_COUT_481_out0;
wire v_COUT_482_out0;
wire v_COUT_483_out0;
wire v_COUT_484_out0;
wire v_COUT_485_out0;
wire v_COUT_486_out0;
wire v_COUT_487_out0;
wire v_COUT_488_out0;
wire v_COUT_489_out0;
wire v_COUT_490_out0;
wire v_COUT_491_out0;
wire v_COUT_492_out0;
wire v_COUT_493_out0;
wire v_COUT_494_out0;
wire v_COUT_495_out0;
wire v_COUT_496_out0;
wire v_COUT_497_out0;
wire v_COUT_498_out0;
wire v_COUT_499_out0;
wire v_COUT_500_out0;
wire v_COUT_501_out0;
wire v_COUT_502_out0;
wire v_COUT_503_out0;
wire v_COUT_504_out0;
wire v_COUT_505_out0;
wire v_COUT_506_out0;
wire v_COUT_507_out0;
wire v_COUT_508_out0;
wire v_COUT_509_out0;
wire v_COUT_510_out0;
wire v_COUT_511_out0;
wire v_COUT_512_out0;
wire v_COUT_513_out0;
wire v_COUT_514_out0;
wire v_COUT_515_out0;
wire v_COUT_516_out0;
wire v_COUT_517_out0;
wire v_COUT_518_out0;
wire v_COUT_5191_out0;
wire v_COUT_519_out0;
wire v_COUT_520_out0;
wire v_COUT_521_out0;
wire v_COUT_522_out0;
wire v_COUT_523_out0;
wire v_COUT_524_out0;
wire v_COUT_525_out0;
wire v_COUT_526_out0;
wire v_COUT_527_out0;
wire v_COUT_528_out0;
wire v_COUT_529_out0;
wire v_COUT_530_out0;
wire v_COUT_531_out0;
wire v_COUT_532_out0;
wire v_COUT_533_out0;
wire v_COUT_534_out0;
wire v_COUT_535_out0;
wire v_COUT_536_out0;
wire v_COUT_537_out0;
wire v_COUT_538_out0;
wire v_COUT_539_out0;
wire v_COUT_540_out0;
wire v_COUT_541_out0;
wire v_COUT_542_out0;
wire v_COUT_543_out0;
wire v_COUT_544_out0;
wire v_COUT_545_out0;
wire v_COUT_546_out0;
wire v_COUT_547_out0;
wire v_COUT_548_out0;
wire v_COUT_549_out0;
wire v_COUT_550_out0;
wire v_COUT_551_out0;
wire v_COUT_552_out0;
wire v_COUT_553_out0;
wire v_COUT_554_out0;
wire v_COUT_555_out0;
wire v_COUT_556_out0;
wire v_C_118_out0;
wire v_C_1559_out0;
wire v_C_1563_out0;
wire v_C_187_out0;
wire v_C_2366_out0;
wire v_C_4256_out0;
wire v_C_4259_out0;
wire v_C_6782_out0;
wire v_D1_4350_out0;
wire v_D1_4350_out1;
wire v_D1_4350_out2;
wire v_D1_4350_out3;
wire v_DIV_INSTRUCTION_1602_out0;
wire v_DIV_INSTRUCTION_2254_out0;
wire v_DIV_INSTRUCTION_5560_out0;
wire v_DIV_INSTRUCTION_6717_out0;
wire v_DONE_RECEIVING_3470_out0;
wire v_D_3773_out0;
wire v_D_3774_out0;
wire v_D_3775_out0;
wire v_D_3776_out0;
wire v_D_3777_out0;
wire v_D_3778_out0;
wire v_D_3779_out0;
wire v_D_3780_out0;
wire v_ENABLE_1292_out0;
wire v_ENABLE_859_out0;
wire v_ENABLE_984_out0;
wire v_ENABLE_985_out0;
wire v_EN_1136_out0;
wire v_EN_1190_out0;
wire v_EN_1423_out0;
wire v_EN_1424_out0;
wire v_EN_1425_out0;
wire v_EN_1426_out0;
wire v_EN_1427_out0;
wire v_EN_1428_out0;
wire v_EN_1429_out0;
wire v_EN_1430_out0;
wire v_EN_2191_out0;
wire v_EN_2243_out0;
wire v_EN_5147_out0;
wire v_EN_5148_out0;
wire v_EN_5158_out0;
wire v_EN_6500_out0;
wire v_EQ01_5173_out0;
wire v_EQ10_1131_out0;
wire v_EQ11_1196_out0;
wire v_EQ1_1238_out0;
wire v_EQ1_1266_out0;
wire v_EQ1_1305_out0;
wire v_EQ1_156_out0;
wire v_EQ1_3415_out0;
wire v_EQ1_3483_out0;
wire v_EQ1_5091_out0;
wire v_EQ1_568_out0;
wire v_EQ1_6617_out0;
wire v_EQ1_907_out0;
wire v_EQ2_3481_out0;
wire v_EQ2_4827_out0;
wire v_EQ2_5099_out0;
wire v_EQ2_5301_out0;
wire v_EQ2_5404_out0;
wire v_EQ2_5540_out0;
wire v_EQ2_5_out0;
wire v_EQ2_6752_out0;
wire v_EQ2_856_out0;
wire v_EQ3_1447_out0;
wire v_EQ3_2871_out0;
wire v_EQ3_3495_out0;
wire v_EQ3_3505_out0;
wire v_EQ3_5434_out0;
wire v_EQ3_6655_out0;
wire v_EQ4_1047_out0;
wire v_EQ4_296_out0;
wire v_EQ4_5098_out0;
wire v_EQ4_560_out0;
wire v_EQ5_2372_out0;
wire v_EQ5_4313_out0;
wire v_EQ5_5106_out0;
wire v_EQ6_11_out0;
wire v_EQ6_827_out0;
wire v_EQ6_961_out0;
wire v_EQ7_1608_out0;
wire v_EQ7_5122_out0;
wire v_EQ8_1194_out0;
wire v_EQ8_1440_out0;
wire v_EQ8_5315_out0;
wire v_EQ9_1165_out0;
wire v_EQ9_2363_out0;
wire v_EQ_1263_out0;
wire v_EQ_1862_out0;
wire v_EQ_52_out0;
wire v_EXEC1LS_209_out0;
wire v_EXEC1LS_2293_out0;
wire v_EXEC1LS_3338_out0;
wire v_EXEC1LS_5171_out0;
wire v_EXEC1LS_5268_out0;
wire v_EXEC1LS_5335_out0;
wire v_EXEC1_1284_out0;
wire v_EXEC1_12_out0;
wire v_EXEC1_1481_out0;
wire v_EXEC1_3451_out0;
wire v_EXEC1_3496_out0;
wire v_EXEC1_5298_out0;
wire v_EXEC1_910_out0;
wire v_EXEC2LS_1389_out0;
wire v_EXEC2LS_1503_out0;
wire v_EXEC2LS_1554_out0;
wire v_EXEC2LS_1573_out0;
wire v_EXEC2LS_5403_out0;
wire v_EXEC2_1290_out0;
wire v_EXEC2_1545_out0;
wire v_EXEC2_1578_out0;
wire v_EXEC2_215_out0;
wire v_EXEC2_3524_out0;
wire v_EXEC2_982_out0;
wire v_EXP1_6644_out0;
wire v_FLAOTING_INSTRUCTION_908_out0;
wire v_FLOATING_EN_ALU_307_out0;
wire v_FLOATING_INSTRUCTION_5118_out0;
wire v_FLOATING_INS_6796_out0;
wire v_FLOAT_2247_out0;
wire v_FLOAT_3772_out0;
wire v_FLOAT_INST16_6621_out0;
wire v_G10_1283_out0;
wire v_G10_1287_out0;
wire v_G10_1288_out0;
wire v_G10_2188_out0;
wire v_G10_292_out0;
wire v_G10_3424_out0;
wire v_G10_3425_out0;
wire v_G10_3426_out0;
wire v_G10_3427_out0;
wire v_G10_3428_out0;
wire v_G10_3429_out0;
wire v_G10_3430_out0;
wire v_G10_3431_out0;
wire v_G10_3432_out0;
wire v_G10_3433_out0;
wire v_G10_3434_out0;
wire v_G10_3435_out0;
wire v_G10_3436_out0;
wire v_G10_3437_out0;
wire v_G10_3438_out0;
wire v_G10_5272_out0;
wire v_G10_6517_out0;
wire v_G10_6518_out0;
wire v_G10_67_out0;
wire v_G10_857_out0;
wire v_G10_950_out0;
wire v_G10_951_out0;
wire v_G11_1243_out0;
wire v_G11_1280_out0;
wire v_G11_1433_out0;
wire v_G11_1434_out0;
wire v_G11_315_out0;
wire v_G11_316_out0;
wire v_G11_317_out0;
wire v_G11_318_out0;
wire v_G11_319_out0;
wire v_G11_320_out0;
wire v_G11_321_out0;
wire v_G11_322_out0;
wire v_G11_323_out0;
wire v_G11_324_out0;
wire v_G11_325_out0;
wire v_G11_326_out0;
wire v_G11_327_out0;
wire v_G11_328_out0;
wire v_G11_329_out0;
wire v_G11_4258_out0;
wire v_G11_5495_out0;
wire v_G11_6572_out0;
wire v_G11_6573_out0;
wire v_G11_6620_out0;
wire v_G12_1107_out0;
wire v_G12_1626_out0;
wire v_G12_1627_out0;
wire v_G12_2294_out0;
wire v_G12_5088_out0;
wire v_G12_5202_out0;
wire v_G12_5261_out0;
wire v_G12_5262_out0;
wire v_G12_6520_out0;
wire v_G12_6521_out0;
wire v_G12_6522_out0;
wire v_G12_6523_out0;
wire v_G12_6524_out0;
wire v_G12_6525_out0;
wire v_G12_6526_out0;
wire v_G12_6527_out0;
wire v_G12_6528_out0;
wire v_G12_6529_out0;
wire v_G12_6530_out0;
wire v_G12_6531_out0;
wire v_G12_6532_out0;
wire v_G12_6533_out0;
wire v_G12_6534_out0;
wire v_G13_2297_out0;
wire v_G13_2298_out0;
wire v_G13_310_out0;
wire v_G13_311_out0;
wire v_G13_3477_out0;
wire v_G13_6577_out0;
wire v_G13_6578_out0;
wire v_G13_6579_out0;
wire v_G13_6580_out0;
wire v_G13_6581_out0;
wire v_G13_6582_out0;
wire v_G13_6583_out0;
wire v_G13_6584_out0;
wire v_G13_6585_out0;
wire v_G13_6586_out0;
wire v_G13_6587_out0;
wire v_G13_6588_out0;
wire v_G13_6589_out0;
wire v_G13_6590_out0;
wire v_G13_6591_out0;
wire v_G14_2215_out0;
wire v_G14_2216_out0;
wire v_G14_298_out0;
wire v_G14_299_out0;
wire v_G14_5126_out0;
wire v_G14_578_out0;
wire v_G14_6542_out0;
wire v_G14_6735_out0;
wire v_G14_6736_out0;
wire v_G14_6737_out0;
wire v_G14_6738_out0;
wire v_G14_6739_out0;
wire v_G14_6740_out0;
wire v_G14_6741_out0;
wire v_G14_6742_out0;
wire v_G14_6743_out0;
wire v_G14_6744_out0;
wire v_G14_6745_out0;
wire v_G14_6746_out0;
wire v_G14_6747_out0;
wire v_G14_6748_out0;
wire v_G14_6749_out0;
wire v_G15_2274_out0;
wire v_G15_2275_out0;
wire v_G15_68_out0;
wire v_G15_69_out0;
wire v_G15_70_out0;
wire v_G15_71_out0;
wire v_G15_72_out0;
wire v_G15_73_out0;
wire v_G15_74_out0;
wire v_G15_75_out0;
wire v_G15_76_out0;
wire v_G15_77_out0;
wire v_G15_78_out0;
wire v_G15_79_out0;
wire v_G15_80_out0;
wire v_G15_81_out0;
wire v_G15_82_out0;
wire v_G15_886_out0;
wire v_G15_887_out0;
wire v_G15_906_out0;
wire v_G16_5365_out0;
wire v_G16_5366_out0;
wire v_G16_5430_out0;
wire v_G16_5431_out0;
wire v_G16_6501_out0;
wire v_G16_6502_out0;
wire v_G16_6503_out0;
wire v_G16_6504_out0;
wire v_G16_6505_out0;
wire v_G16_6506_out0;
wire v_G16_6507_out0;
wire v_G16_6508_out0;
wire v_G16_6509_out0;
wire v_G16_6510_out0;
wire v_G16_6511_out0;
wire v_G16_6512_out0;
wire v_G16_6513_out0;
wire v_G16_6514_out0;
wire v_G16_6515_out0;
wire v_G16_6595_out0;
wire v_G18_4330_out0;
wire v_G18_4331_out0;
wire v_G18_5514_out0;
wire v_G19_2277_out0;
wire v_G1_1085_out0;
wire v_G1_1318_out0;
wire v_G1_1319_out0;
wire v_G1_1320_out0;
wire v_G1_1321_out0;
wire v_G1_1322_out0;
wire v_G1_1323_out0;
wire v_G1_1324_out0;
wire v_G1_1325_out0;
wire v_G1_138_out0;
wire v_G1_1418_out0;
wire v_G1_143_out0;
wire v_G1_1473_out0;
wire v_G1_1949_out0;
wire v_G1_1950_out0;
wire v_G1_1951_out0;
wire v_G1_1952_out0;
wire v_G1_1953_out0;
wire v_G1_1954_out0;
wire v_G1_1955_out0;
wire v_G1_1956_out0;
wire v_G1_1957_out0;
wire v_G1_1958_out0;
wire v_G1_1959_out0;
wire v_G1_1960_out0;
wire v_G1_1961_out0;
wire v_G1_1962_out0;
wire v_G1_1963_out0;
wire v_G1_1964_out0;
wire v_G1_1965_out0;
wire v_G1_1966_out0;
wire v_G1_1967_out0;
wire v_G1_1968_out0;
wire v_G1_1969_out0;
wire v_G1_1970_out0;
wire v_G1_1971_out0;
wire v_G1_1972_out0;
wire v_G1_1973_out0;
wire v_G1_1974_out0;
wire v_G1_1975_out0;
wire v_G1_1976_out0;
wire v_G1_1977_out0;
wire v_G1_1978_out0;
wire v_G1_1979_out0;
wire v_G1_1980_out0;
wire v_G1_1981_out0;
wire v_G1_1982_out0;
wire v_G1_1983_out0;
wire v_G1_1984_out0;
wire v_G1_1985_out0;
wire v_G1_1986_out0;
wire v_G1_1987_out0;
wire v_G1_1988_out0;
wire v_G1_1989_out0;
wire v_G1_1990_out0;
wire v_G1_1991_out0;
wire v_G1_1992_out0;
wire v_G1_1993_out0;
wire v_G1_1994_out0;
wire v_G1_1995_out0;
wire v_G1_1996_out0;
wire v_G1_1997_out0;
wire v_G1_1998_out0;
wire v_G1_1999_out0;
wire v_G1_2000_out0;
wire v_G1_2001_out0;
wire v_G1_2002_out0;
wire v_G1_2003_out0;
wire v_G1_2004_out0;
wire v_G1_2005_out0;
wire v_G1_2006_out0;
wire v_G1_2007_out0;
wire v_G1_2008_out0;
wire v_G1_2009_out0;
wire v_G1_2010_out0;
wire v_G1_2011_out0;
wire v_G1_2012_out0;
wire v_G1_2013_out0;
wire v_G1_2014_out0;
wire v_G1_2015_out0;
wire v_G1_2016_out0;
wire v_G1_2017_out0;
wire v_G1_2018_out0;
wire v_G1_2019_out0;
wire v_G1_2020_out0;
wire v_G1_2021_out0;
wire v_G1_2022_out0;
wire v_G1_2023_out0;
wire v_G1_2024_out0;
wire v_G1_2025_out0;
wire v_G1_2026_out0;
wire v_G1_2027_out0;
wire v_G1_2028_out0;
wire v_G1_2029_out0;
wire v_G1_2030_out0;
wire v_G1_2031_out0;
wire v_G1_2032_out0;
wire v_G1_2033_out0;
wire v_G1_2034_out0;
wire v_G1_2035_out0;
wire v_G1_2036_out0;
wire v_G1_2037_out0;
wire v_G1_2038_out0;
wire v_G1_2039_out0;
wire v_G1_2040_out0;
wire v_G1_2041_out0;
wire v_G1_2042_out0;
wire v_G1_2043_out0;
wire v_G1_2044_out0;
wire v_G1_2045_out0;
wire v_G1_2046_out0;
wire v_G1_2047_out0;
wire v_G1_2048_out0;
wire v_G1_2049_out0;
wire v_G1_2050_out0;
wire v_G1_2051_out0;
wire v_G1_2052_out0;
wire v_G1_2053_out0;
wire v_G1_2054_out0;
wire v_G1_2055_out0;
wire v_G1_2056_out0;
wire v_G1_2057_out0;
wire v_G1_2058_out0;
wire v_G1_2059_out0;
wire v_G1_2060_out0;
wire v_G1_2061_out0;
wire v_G1_2062_out0;
wire v_G1_2063_out0;
wire v_G1_2064_out0;
wire v_G1_2065_out0;
wire v_G1_2066_out0;
wire v_G1_2067_out0;
wire v_G1_2068_out0;
wire v_G1_2069_out0;
wire v_G1_2070_out0;
wire v_G1_2071_out0;
wire v_G1_2072_out0;
wire v_G1_2073_out0;
wire v_G1_2074_out0;
wire v_G1_2075_out0;
wire v_G1_2076_out0;
wire v_G1_2077_out0;
wire v_G1_2078_out0;
wire v_G1_2079_out0;
wire v_G1_2080_out0;
wire v_G1_2081_out0;
wire v_G1_2082_out0;
wire v_G1_2083_out0;
wire v_G1_2084_out0;
wire v_G1_2085_out0;
wire v_G1_2086_out0;
wire v_G1_2087_out0;
wire v_G1_2088_out0;
wire v_G1_2089_out0;
wire v_G1_2090_out0;
wire v_G1_2091_out0;
wire v_G1_2092_out0;
wire v_G1_2093_out0;
wire v_G1_2094_out0;
wire v_G1_2095_out0;
wire v_G1_2096_out0;
wire v_G1_2097_out0;
wire v_G1_2098_out0;
wire v_G1_2099_out0;
wire v_G1_2100_out0;
wire v_G1_2101_out0;
wire v_G1_2102_out0;
wire v_G1_2103_out0;
wire v_G1_2104_out0;
wire v_G1_2105_out0;
wire v_G1_2106_out0;
wire v_G1_2107_out0;
wire v_G1_2108_out0;
wire v_G1_2109_out0;
wire v_G1_2110_out0;
wire v_G1_2111_out0;
wire v_G1_2112_out0;
wire v_G1_2113_out0;
wire v_G1_2114_out0;
wire v_G1_2115_out0;
wire v_G1_2116_out0;
wire v_G1_2117_out0;
wire v_G1_2118_out0;
wire v_G1_2119_out0;
wire v_G1_2120_out0;
wire v_G1_2121_out0;
wire v_G1_2122_out0;
wire v_G1_2123_out0;
wire v_G1_2124_out0;
wire v_G1_2125_out0;
wire v_G1_2126_out0;
wire v_G1_2127_out0;
wire v_G1_2128_out0;
wire v_G1_2129_out0;
wire v_G1_2130_out0;
wire v_G1_2131_out0;
wire v_G1_2132_out0;
wire v_G1_2133_out0;
wire v_G1_2134_out0;
wire v_G1_2135_out0;
wire v_G1_2136_out0;
wire v_G1_2137_out0;
wire v_G1_2138_out0;
wire v_G1_2139_out0;
wire v_G1_2140_out0;
wire v_G1_2141_out0;
wire v_G1_2142_out0;
wire v_G1_2143_out0;
wire v_G1_2144_out0;
wire v_G1_2145_out0;
wire v_G1_2146_out0;
wire v_G1_2147_out0;
wire v_G1_2148_out0;
wire v_G1_2149_out0;
wire v_G1_2150_out0;
wire v_G1_2151_out0;
wire v_G1_2152_out0;
wire v_G1_2153_out0;
wire v_G1_2154_out0;
wire v_G1_2155_out0;
wire v_G1_2156_out0;
wire v_G1_2157_out0;
wire v_G1_2158_out0;
wire v_G1_2159_out0;
wire v_G1_2160_out0;
wire v_G1_2161_out0;
wire v_G1_2162_out0;
wire v_G1_2163_out0;
wire v_G1_2164_out0;
wire v_G1_2165_out0;
wire v_G1_2166_out0;
wire v_G1_2167_out0;
wire v_G1_2168_out0;
wire v_G1_2169_out0;
wire v_G1_2170_out0;
wire v_G1_2171_out0;
wire v_G1_2172_out0;
wire v_G1_312_out0;
wire v_G1_3791_out0;
wire v_G1_3792_out0;
wire v_G1_3793_out0;
wire v_G1_3794_out0;
wire v_G1_3795_out0;
wire v_G1_3796_out0;
wire v_G1_3797_out0;
wire v_G1_3798_out0;
wire v_G1_3799_out0;
wire v_G1_3800_out0;
wire v_G1_3801_out0;
wire v_G1_3802_out0;
wire v_G1_3803_out0;
wire v_G1_3804_out0;
wire v_G1_3805_out0;
wire v_G1_3806_out0;
wire v_G1_3807_out0;
wire v_G1_3808_out0;
wire v_G1_3809_out0;
wire v_G1_3810_out0;
wire v_G1_3811_out0;
wire v_G1_3812_out0;
wire v_G1_3813_out0;
wire v_G1_3814_out0;
wire v_G1_3815_out0;
wire v_G1_3816_out0;
wire v_G1_3817_out0;
wire v_G1_3818_out0;
wire v_G1_3819_out0;
wire v_G1_3820_out0;
wire v_G1_3821_out0;
wire v_G1_3822_out0;
wire v_G1_3823_out0;
wire v_G1_3824_out0;
wire v_G1_3825_out0;
wire v_G1_3826_out0;
wire v_G1_3827_out0;
wire v_G1_3828_out0;
wire v_G1_3829_out0;
wire v_G1_3830_out0;
wire v_G1_3831_out0;
wire v_G1_3832_out0;
wire v_G1_3833_out0;
wire v_G1_3834_out0;
wire v_G1_3835_out0;
wire v_G1_3836_out0;
wire v_G1_3837_out0;
wire v_G1_3838_out0;
wire v_G1_3839_out0;
wire v_G1_3840_out0;
wire v_G1_3841_out0;
wire v_G1_3842_out0;
wire v_G1_3843_out0;
wire v_G1_3844_out0;
wire v_G1_3845_out0;
wire v_G1_3846_out0;
wire v_G1_3847_out0;
wire v_G1_3848_out0;
wire v_G1_3849_out0;
wire v_G1_3850_out0;
wire v_G1_3851_out0;
wire v_G1_3852_out0;
wire v_G1_3853_out0;
wire v_G1_3854_out0;
wire v_G1_3855_out0;
wire v_G1_3856_out0;
wire v_G1_3857_out0;
wire v_G1_3858_out0;
wire v_G1_3859_out0;
wire v_G1_3860_out0;
wire v_G1_3861_out0;
wire v_G1_3862_out0;
wire v_G1_3863_out0;
wire v_G1_3864_out0;
wire v_G1_3865_out0;
wire v_G1_3866_out0;
wire v_G1_3867_out0;
wire v_G1_3868_out0;
wire v_G1_3869_out0;
wire v_G1_3870_out0;
wire v_G1_3871_out0;
wire v_G1_3872_out0;
wire v_G1_3873_out0;
wire v_G1_3874_out0;
wire v_G1_3875_out0;
wire v_G1_3876_out0;
wire v_G1_3877_out0;
wire v_G1_3878_out0;
wire v_G1_3879_out0;
wire v_G1_3880_out0;
wire v_G1_3881_out0;
wire v_G1_3882_out0;
wire v_G1_3883_out0;
wire v_G1_3884_out0;
wire v_G1_3885_out0;
wire v_G1_3886_out0;
wire v_G1_3887_out0;
wire v_G1_3888_out0;
wire v_G1_3889_out0;
wire v_G1_3890_out0;
wire v_G1_3891_out0;
wire v_G1_3892_out0;
wire v_G1_3893_out0;
wire v_G1_3894_out0;
wire v_G1_3895_out0;
wire v_G1_3896_out0;
wire v_G1_3897_out0;
wire v_G1_3898_out0;
wire v_G1_3899_out0;
wire v_G1_3900_out0;
wire v_G1_3901_out0;
wire v_G1_3902_out0;
wire v_G1_3903_out0;
wire v_G1_3904_out0;
wire v_G1_3905_out0;
wire v_G1_3906_out0;
wire v_G1_3907_out0;
wire v_G1_3908_out0;
wire v_G1_3909_out0;
wire v_G1_3910_out0;
wire v_G1_3911_out0;
wire v_G1_3912_out0;
wire v_G1_3913_out0;
wire v_G1_3914_out0;
wire v_G1_3915_out0;
wire v_G1_3916_out0;
wire v_G1_3917_out0;
wire v_G1_3918_out0;
wire v_G1_3919_out0;
wire v_G1_3920_out0;
wire v_G1_3921_out0;
wire v_G1_3922_out0;
wire v_G1_3923_out0;
wire v_G1_3924_out0;
wire v_G1_3925_out0;
wire v_G1_3926_out0;
wire v_G1_3927_out0;
wire v_G1_3928_out0;
wire v_G1_3929_out0;
wire v_G1_3930_out0;
wire v_G1_3931_out0;
wire v_G1_3932_out0;
wire v_G1_3933_out0;
wire v_G1_3934_out0;
wire v_G1_3935_out0;
wire v_G1_3936_out0;
wire v_G1_3937_out0;
wire v_G1_3938_out0;
wire v_G1_3939_out0;
wire v_G1_3940_out0;
wire v_G1_3941_out0;
wire v_G1_3942_out0;
wire v_G1_3943_out0;
wire v_G1_3944_out0;
wire v_G1_3945_out0;
wire v_G1_3946_out0;
wire v_G1_3947_out0;
wire v_G1_3948_out0;
wire v_G1_3949_out0;
wire v_G1_3950_out0;
wire v_G1_3951_out0;
wire v_G1_3952_out0;
wire v_G1_3953_out0;
wire v_G1_3954_out0;
wire v_G1_3955_out0;
wire v_G1_3956_out0;
wire v_G1_3957_out0;
wire v_G1_3958_out0;
wire v_G1_3959_out0;
wire v_G1_3960_out0;
wire v_G1_3961_out0;
wire v_G1_3962_out0;
wire v_G1_3963_out0;
wire v_G1_3964_out0;
wire v_G1_3965_out0;
wire v_G1_3966_out0;
wire v_G1_3967_out0;
wire v_G1_3968_out0;
wire v_G1_3969_out0;
wire v_G1_3970_out0;
wire v_G1_3971_out0;
wire v_G1_3972_out0;
wire v_G1_3973_out0;
wire v_G1_3974_out0;
wire v_G1_3975_out0;
wire v_G1_3976_out0;
wire v_G1_3977_out0;
wire v_G1_3978_out0;
wire v_G1_3979_out0;
wire v_G1_3980_out0;
wire v_G1_3981_out0;
wire v_G1_3982_out0;
wire v_G1_3983_out0;
wire v_G1_3984_out0;
wire v_G1_3985_out0;
wire v_G1_3986_out0;
wire v_G1_3987_out0;
wire v_G1_3988_out0;
wire v_G1_3989_out0;
wire v_G1_3990_out0;
wire v_G1_3991_out0;
wire v_G1_3992_out0;
wire v_G1_3993_out0;
wire v_G1_3994_out0;
wire v_G1_3995_out0;
wire v_G1_3996_out0;
wire v_G1_3997_out0;
wire v_G1_3998_out0;
wire v_G1_3999_out0;
wire v_G1_4000_out0;
wire v_G1_4001_out0;
wire v_G1_4002_out0;
wire v_G1_4003_out0;
wire v_G1_4004_out0;
wire v_G1_4005_out0;
wire v_G1_4006_out0;
wire v_G1_4007_out0;
wire v_G1_4008_out0;
wire v_G1_4009_out0;
wire v_G1_4010_out0;
wire v_G1_4011_out0;
wire v_G1_4012_out0;
wire v_G1_4013_out0;
wire v_G1_4014_out0;
wire v_G1_4015_out0;
wire v_G1_4016_out0;
wire v_G1_4017_out0;
wire v_G1_4018_out0;
wire v_G1_4019_out0;
wire v_G1_4020_out0;
wire v_G1_4021_out0;
wire v_G1_4022_out0;
wire v_G1_4023_out0;
wire v_G1_4024_out0;
wire v_G1_4025_out0;
wire v_G1_4026_out0;
wire v_G1_4027_out0;
wire v_G1_4028_out0;
wire v_G1_4029_out0;
wire v_G1_4030_out0;
wire v_G1_4031_out0;
wire v_G1_4032_out0;
wire v_G1_4033_out0;
wire v_G1_4034_out0;
wire v_G1_4035_out0;
wire v_G1_4036_out0;
wire v_G1_4037_out0;
wire v_G1_4038_out0;
wire v_G1_4039_out0;
wire v_G1_4040_out0;
wire v_G1_4041_out0;
wire v_G1_4042_out0;
wire v_G1_4043_out0;
wire v_G1_4044_out0;
wire v_G1_4045_out0;
wire v_G1_4046_out0;
wire v_G1_4047_out0;
wire v_G1_4048_out0;
wire v_G1_4049_out0;
wire v_G1_4050_out0;
wire v_G1_4051_out0;
wire v_G1_4052_out0;
wire v_G1_4053_out0;
wire v_G1_4054_out0;
wire v_G1_4055_out0;
wire v_G1_4056_out0;
wire v_G1_4057_out0;
wire v_G1_4058_out0;
wire v_G1_4059_out0;
wire v_G1_4060_out0;
wire v_G1_4061_out0;
wire v_G1_4062_out0;
wire v_G1_4063_out0;
wire v_G1_4064_out0;
wire v_G1_4065_out0;
wire v_G1_4066_out0;
wire v_G1_4067_out0;
wire v_G1_4068_out0;
wire v_G1_4069_out0;
wire v_G1_4070_out0;
wire v_G1_4071_out0;
wire v_G1_4072_out0;
wire v_G1_4073_out0;
wire v_G1_4074_out0;
wire v_G1_4075_out0;
wire v_G1_4076_out0;
wire v_G1_4077_out0;
wire v_G1_4078_out0;
wire v_G1_4079_out0;
wire v_G1_4080_out0;
wire v_G1_4081_out0;
wire v_G1_4082_out0;
wire v_G1_4083_out0;
wire v_G1_4084_out0;
wire v_G1_4085_out0;
wire v_G1_4086_out0;
wire v_G1_4087_out0;
wire v_G1_4088_out0;
wire v_G1_4089_out0;
wire v_G1_4090_out0;
wire v_G1_4091_out0;
wire v_G1_4092_out0;
wire v_G1_4093_out0;
wire v_G1_4094_out0;
wire v_G1_4095_out0;
wire v_G1_4096_out0;
wire v_G1_4097_out0;
wire v_G1_4098_out0;
wire v_G1_4099_out0;
wire v_G1_4100_out0;
wire v_G1_4101_out0;
wire v_G1_4102_out0;
wire v_G1_4103_out0;
wire v_G1_4104_out0;
wire v_G1_4105_out0;
wire v_G1_4106_out0;
wire v_G1_4107_out0;
wire v_G1_4108_out0;
wire v_G1_4109_out0;
wire v_G1_4110_out0;
wire v_G1_4111_out0;
wire v_G1_4112_out0;
wire v_G1_4113_out0;
wire v_G1_4114_out0;
wire v_G1_4115_out0;
wire v_G1_4116_out0;
wire v_G1_4117_out0;
wire v_G1_4118_out0;
wire v_G1_4119_out0;
wire v_G1_4120_out0;
wire v_G1_4121_out0;
wire v_G1_4122_out0;
wire v_G1_4123_out0;
wire v_G1_4124_out0;
wire v_G1_4125_out0;
wire v_G1_4126_out0;
wire v_G1_4127_out0;
wire v_G1_4128_out0;
wire v_G1_4129_out0;
wire v_G1_4130_out0;
wire v_G1_4131_out0;
wire v_G1_4132_out0;
wire v_G1_4133_out0;
wire v_G1_4134_out0;
wire v_G1_4135_out0;
wire v_G1_4136_out0;
wire v_G1_4137_out0;
wire v_G1_4138_out0;
wire v_G1_4139_out0;
wire v_G1_4140_out0;
wire v_G1_4141_out0;
wire v_G1_4142_out0;
wire v_G1_4143_out0;
wire v_G1_4144_out0;
wire v_G1_4145_out0;
wire v_G1_4146_out0;
wire v_G1_4147_out0;
wire v_G1_4148_out0;
wire v_G1_4149_out0;
wire v_G1_4150_out0;
wire v_G1_4151_out0;
wire v_G1_4152_out0;
wire v_G1_4153_out0;
wire v_G1_4154_out0;
wire v_G1_4155_out0;
wire v_G1_4156_out0;
wire v_G1_4157_out0;
wire v_G1_4158_out0;
wire v_G1_4159_out0;
wire v_G1_4160_out0;
wire v_G1_4161_out0;
wire v_G1_4162_out0;
wire v_G1_4163_out0;
wire v_G1_4164_out0;
wire v_G1_4165_out0;
wire v_G1_4166_out0;
wire v_G1_4167_out0;
wire v_G1_4168_out0;
wire v_G1_4169_out0;
wire v_G1_4170_out0;
wire v_G1_4171_out0;
wire v_G1_4172_out0;
wire v_G1_4173_out0;
wire v_G1_4174_out0;
wire v_G1_4175_out0;
wire v_G1_4176_out0;
wire v_G1_4177_out0;
wire v_G1_4178_out0;
wire v_G1_4179_out0;
wire v_G1_4180_out0;
wire v_G1_4181_out0;
wire v_G1_4182_out0;
wire v_G1_4183_out0;
wire v_G1_4184_out0;
wire v_G1_4185_out0;
wire v_G1_4186_out0;
wire v_G1_4187_out0;
wire v_G1_4188_out0;
wire v_G1_4189_out0;
wire v_G1_4190_out0;
wire v_G1_4191_out0;
wire v_G1_4192_out0;
wire v_G1_4193_out0;
wire v_G1_4194_out0;
wire v_G1_4195_out0;
wire v_G1_4196_out0;
wire v_G1_4197_out0;
wire v_G1_4198_out0;
wire v_G1_4199_out0;
wire v_G1_4200_out0;
wire v_G1_4201_out0;
wire v_G1_4202_out0;
wire v_G1_4203_out0;
wire v_G1_4204_out0;
wire v_G1_4205_out0;
wire v_G1_4206_out0;
wire v_G1_4207_out0;
wire v_G1_4208_out0;
wire v_G1_4209_out0;
wire v_G1_4210_out0;
wire v_G1_4211_out0;
wire v_G1_4212_out0;
wire v_G1_4213_out0;
wire v_G1_4214_out0;
wire v_G1_4215_out0;
wire v_G1_4216_out0;
wire v_G1_4217_out0;
wire v_G1_4218_out0;
wire v_G1_4219_out0;
wire v_G1_4220_out0;
wire v_G1_4221_out0;
wire v_G1_4222_out0;
wire v_G1_4223_out0;
wire v_G1_4224_out0;
wire v_G1_4225_out0;
wire v_G1_4226_out0;
wire v_G1_4227_out0;
wire v_G1_4228_out0;
wire v_G1_4229_out0;
wire v_G1_4230_out0;
wire v_G1_4231_out0;
wire v_G1_4232_out0;
wire v_G1_4233_out0;
wire v_G1_4234_out0;
wire v_G1_4235_out0;
wire v_G1_4236_out0;
wire v_G1_4237_out0;
wire v_G1_4238_out0;
wire v_G1_4239_out0;
wire v_G1_4240_out0;
wire v_G1_4241_out0;
wire v_G1_4242_out0;
wire v_G1_4243_out0;
wire v_G1_4244_out0;
wire v_G1_4245_out0;
wire v_G1_4246_out0;
wire v_G1_4247_out0;
wire v_G1_4248_out0;
wire v_G1_4249_out0;
wire v_G1_4250_out0;
wire v_G1_4251_out0;
wire v_G1_4252_out0;
wire v_G1_4253_out0;
wire v_G1_4254_out0;
wire v_G1_4279_out0;
wire v_G1_4280_out0;
wire v_G1_5159_out0;
wire v_G1_5271_out0;
wire v_G1_5295_out0;
wire v_G1_5318_out0;
wire v_G1_5491_out0;
wire v_G1_573_out0;
wire v_G1_583_out0;
wire v_G1_6776_out0;
wire v_G1_6777_out0;
wire v_G1_6786_out0;
wire v_G1_919_out0;
wire v_G1_920_out0;
wire v_G1_933_out0;
wire v_G1_934_out0;
wire v_G1_935_out0;
wire v_G1_936_out0;
wire v_G1_937_out0;
wire v_G1_938_out0;
wire v_G1_939_out0;
wire v_G1_940_out0;
wire v_G1_941_out0;
wire v_G1_942_out0;
wire v_G1_943_out0;
wire v_G1_944_out0;
wire v_G1_945_out0;
wire v_G1_946_out0;
wire v_G1_947_out0;
wire v_G20_5486_out0;
wire v_G21_1405_out0;
wire v_G21_1856_out0;
wire v_G21_1857_out0;
wire v_G22_5405_out0;
wire v_G22_5406_out0;
wire v_G23_1387_out0;
wire v_G23_2368_out0;
wire v_G23_2369_out0;
wire v_G24_1930_out0;
wire v_G24_5196_out0;
wire v_G24_5197_out0;
wire v_G25_3418_out0;
wire v_G26_2312_out0;
wire v_G27_4825_out0;
wire v_G28_1025_out0;
wire v_G28_1026_out0;
wire v_G28_3373_out0;
wire v_G29_2860_out0;
wire v_G2_1293_out0;
wire v_G2_1408_out0;
wire v_G2_1452_out0;
wire v_G2_1453_out0;
wire v_G2_1569_out0;
wire v_G2_1577_out0;
wire v_G2_1579_out0;
wire v_G2_2257_out0;
wire v_G2_2258_out0;
wire v_G2_2259_out0;
wire v_G2_2260_out0;
wire v_G2_2261_out0;
wire v_G2_2262_out0;
wire v_G2_2263_out0;
wire v_G2_2264_out0;
wire v_G2_2265_out0;
wire v_G2_2266_out0;
wire v_G2_2267_out0;
wire v_G2_2268_out0;
wire v_G2_2269_out0;
wire v_G2_2270_out0;
wire v_G2_2271_out0;
wire v_G2_2863_out0;
wire v_G2_3336_out0;
wire v_G2_3380_out0;
wire v_G2_3444_out0;
wire v_G2_3449_out0;
wire v_G2_3450_out0;
wire v_G2_5068_out0;
wire v_G2_5156_out0;
wire v_G2_5313_out0;
wire v_G2_5481_out0;
wire v_G2_6027_out0;
wire v_G2_6036_out0;
wire v_G2_6037_out0;
wire v_G2_6038_out0;
wire v_G2_6039_out0;
wire v_G2_6040_out0;
wire v_G2_6041_out0;
wire v_G2_6042_out0;
wire v_G2_6043_out0;
wire v_G2_6044_out0;
wire v_G2_6045_out0;
wire v_G2_6046_out0;
wire v_G2_6047_out0;
wire v_G2_6048_out0;
wire v_G2_6049_out0;
wire v_G2_6050_out0;
wire v_G2_6051_out0;
wire v_G2_6052_out0;
wire v_G2_6053_out0;
wire v_G2_6054_out0;
wire v_G2_6055_out0;
wire v_G2_6056_out0;
wire v_G2_6057_out0;
wire v_G2_6058_out0;
wire v_G2_6059_out0;
wire v_G2_6060_out0;
wire v_G2_6061_out0;
wire v_G2_6062_out0;
wire v_G2_6063_out0;
wire v_G2_6064_out0;
wire v_G2_6065_out0;
wire v_G2_6066_out0;
wire v_G2_6067_out0;
wire v_G2_6068_out0;
wire v_G2_6069_out0;
wire v_G2_6070_out0;
wire v_G2_6071_out0;
wire v_G2_6072_out0;
wire v_G2_6073_out0;
wire v_G2_6074_out0;
wire v_G2_6075_out0;
wire v_G2_6076_out0;
wire v_G2_6077_out0;
wire v_G2_6078_out0;
wire v_G2_6079_out0;
wire v_G2_6080_out0;
wire v_G2_6081_out0;
wire v_G2_6082_out0;
wire v_G2_6083_out0;
wire v_G2_6084_out0;
wire v_G2_6085_out0;
wire v_G2_6086_out0;
wire v_G2_6087_out0;
wire v_G2_6088_out0;
wire v_G2_6089_out0;
wire v_G2_6090_out0;
wire v_G2_6091_out0;
wire v_G2_6092_out0;
wire v_G2_6093_out0;
wire v_G2_6094_out0;
wire v_G2_6095_out0;
wire v_G2_6096_out0;
wire v_G2_6097_out0;
wire v_G2_6098_out0;
wire v_G2_6099_out0;
wire v_G2_6100_out0;
wire v_G2_6101_out0;
wire v_G2_6102_out0;
wire v_G2_6103_out0;
wire v_G2_6104_out0;
wire v_G2_6105_out0;
wire v_G2_6106_out0;
wire v_G2_6107_out0;
wire v_G2_6108_out0;
wire v_G2_6109_out0;
wire v_G2_6110_out0;
wire v_G2_6111_out0;
wire v_G2_6112_out0;
wire v_G2_6113_out0;
wire v_G2_6114_out0;
wire v_G2_6115_out0;
wire v_G2_6116_out0;
wire v_G2_6117_out0;
wire v_G2_6118_out0;
wire v_G2_6119_out0;
wire v_G2_6120_out0;
wire v_G2_6121_out0;
wire v_G2_6122_out0;
wire v_G2_6123_out0;
wire v_G2_6124_out0;
wire v_G2_6125_out0;
wire v_G2_6126_out0;
wire v_G2_6127_out0;
wire v_G2_6128_out0;
wire v_G2_6129_out0;
wire v_G2_6130_out0;
wire v_G2_6131_out0;
wire v_G2_6132_out0;
wire v_G2_6133_out0;
wire v_G2_6134_out0;
wire v_G2_6135_out0;
wire v_G2_6136_out0;
wire v_G2_6137_out0;
wire v_G2_6138_out0;
wire v_G2_6139_out0;
wire v_G2_6140_out0;
wire v_G2_6141_out0;
wire v_G2_6142_out0;
wire v_G2_6143_out0;
wire v_G2_6144_out0;
wire v_G2_6145_out0;
wire v_G2_6146_out0;
wire v_G2_6147_out0;
wire v_G2_6148_out0;
wire v_G2_6149_out0;
wire v_G2_6150_out0;
wire v_G2_6151_out0;
wire v_G2_6152_out0;
wire v_G2_6153_out0;
wire v_G2_6154_out0;
wire v_G2_6155_out0;
wire v_G2_6156_out0;
wire v_G2_6157_out0;
wire v_G2_6158_out0;
wire v_G2_6159_out0;
wire v_G2_6160_out0;
wire v_G2_6161_out0;
wire v_G2_6162_out0;
wire v_G2_6163_out0;
wire v_G2_6164_out0;
wire v_G2_6165_out0;
wire v_G2_6166_out0;
wire v_G2_6167_out0;
wire v_G2_6168_out0;
wire v_G2_6169_out0;
wire v_G2_6170_out0;
wire v_G2_6171_out0;
wire v_G2_6172_out0;
wire v_G2_6173_out0;
wire v_G2_6174_out0;
wire v_G2_6175_out0;
wire v_G2_6176_out0;
wire v_G2_6177_out0;
wire v_G2_6178_out0;
wire v_G2_6179_out0;
wire v_G2_6180_out0;
wire v_G2_6181_out0;
wire v_G2_6182_out0;
wire v_G2_6183_out0;
wire v_G2_6184_out0;
wire v_G2_6185_out0;
wire v_G2_6186_out0;
wire v_G2_6187_out0;
wire v_G2_6188_out0;
wire v_G2_6189_out0;
wire v_G2_6190_out0;
wire v_G2_6191_out0;
wire v_G2_6192_out0;
wire v_G2_6193_out0;
wire v_G2_6194_out0;
wire v_G2_6195_out0;
wire v_G2_6196_out0;
wire v_G2_6197_out0;
wire v_G2_6198_out0;
wire v_G2_6199_out0;
wire v_G2_6200_out0;
wire v_G2_6201_out0;
wire v_G2_6202_out0;
wire v_G2_6203_out0;
wire v_G2_6204_out0;
wire v_G2_6205_out0;
wire v_G2_6206_out0;
wire v_G2_6207_out0;
wire v_G2_6208_out0;
wire v_G2_6209_out0;
wire v_G2_6210_out0;
wire v_G2_6211_out0;
wire v_G2_6212_out0;
wire v_G2_6213_out0;
wire v_G2_6214_out0;
wire v_G2_6215_out0;
wire v_G2_6216_out0;
wire v_G2_6217_out0;
wire v_G2_6218_out0;
wire v_G2_6219_out0;
wire v_G2_6220_out0;
wire v_G2_6221_out0;
wire v_G2_6222_out0;
wire v_G2_6223_out0;
wire v_G2_6224_out0;
wire v_G2_6225_out0;
wire v_G2_6226_out0;
wire v_G2_6227_out0;
wire v_G2_6228_out0;
wire v_G2_6229_out0;
wire v_G2_6230_out0;
wire v_G2_6231_out0;
wire v_G2_6232_out0;
wire v_G2_6233_out0;
wire v_G2_6234_out0;
wire v_G2_6235_out0;
wire v_G2_6236_out0;
wire v_G2_6237_out0;
wire v_G2_6238_out0;
wire v_G2_6239_out0;
wire v_G2_6240_out0;
wire v_G2_6241_out0;
wire v_G2_6242_out0;
wire v_G2_6243_out0;
wire v_G2_6244_out0;
wire v_G2_6245_out0;
wire v_G2_6246_out0;
wire v_G2_6247_out0;
wire v_G2_6248_out0;
wire v_G2_6249_out0;
wire v_G2_6250_out0;
wire v_G2_6251_out0;
wire v_G2_6252_out0;
wire v_G2_6253_out0;
wire v_G2_6254_out0;
wire v_G2_6255_out0;
wire v_G2_6256_out0;
wire v_G2_6257_out0;
wire v_G2_6258_out0;
wire v_G2_6259_out0;
wire v_G2_6260_out0;
wire v_G2_6261_out0;
wire v_G2_6262_out0;
wire v_G2_6263_out0;
wire v_G2_6264_out0;
wire v_G2_6265_out0;
wire v_G2_6266_out0;
wire v_G2_6267_out0;
wire v_G2_6268_out0;
wire v_G2_6269_out0;
wire v_G2_6270_out0;
wire v_G2_6271_out0;
wire v_G2_6272_out0;
wire v_G2_6273_out0;
wire v_G2_6274_out0;
wire v_G2_6275_out0;
wire v_G2_6276_out0;
wire v_G2_6277_out0;
wire v_G2_6278_out0;
wire v_G2_6279_out0;
wire v_G2_6280_out0;
wire v_G2_6281_out0;
wire v_G2_6282_out0;
wire v_G2_6283_out0;
wire v_G2_6284_out0;
wire v_G2_6285_out0;
wire v_G2_6286_out0;
wire v_G2_6287_out0;
wire v_G2_6288_out0;
wire v_G2_6289_out0;
wire v_G2_6290_out0;
wire v_G2_6291_out0;
wire v_G2_6292_out0;
wire v_G2_6293_out0;
wire v_G2_6294_out0;
wire v_G2_6295_out0;
wire v_G2_6296_out0;
wire v_G2_6297_out0;
wire v_G2_6298_out0;
wire v_G2_6299_out0;
wire v_G2_6300_out0;
wire v_G2_6301_out0;
wire v_G2_6302_out0;
wire v_G2_6303_out0;
wire v_G2_6304_out0;
wire v_G2_6305_out0;
wire v_G2_6306_out0;
wire v_G2_6307_out0;
wire v_G2_6308_out0;
wire v_G2_6309_out0;
wire v_G2_6310_out0;
wire v_G2_6311_out0;
wire v_G2_6312_out0;
wire v_G2_6313_out0;
wire v_G2_6314_out0;
wire v_G2_6315_out0;
wire v_G2_6316_out0;
wire v_G2_6317_out0;
wire v_G2_6318_out0;
wire v_G2_6319_out0;
wire v_G2_6320_out0;
wire v_G2_6321_out0;
wire v_G2_6322_out0;
wire v_G2_6323_out0;
wire v_G2_6324_out0;
wire v_G2_6325_out0;
wire v_G2_6326_out0;
wire v_G2_6327_out0;
wire v_G2_6328_out0;
wire v_G2_6329_out0;
wire v_G2_6330_out0;
wire v_G2_6331_out0;
wire v_G2_6332_out0;
wire v_G2_6333_out0;
wire v_G2_6334_out0;
wire v_G2_6335_out0;
wire v_G2_6336_out0;
wire v_G2_6337_out0;
wire v_G2_6338_out0;
wire v_G2_6339_out0;
wire v_G2_6340_out0;
wire v_G2_6341_out0;
wire v_G2_6342_out0;
wire v_G2_6343_out0;
wire v_G2_6344_out0;
wire v_G2_6345_out0;
wire v_G2_6346_out0;
wire v_G2_6347_out0;
wire v_G2_6348_out0;
wire v_G2_6349_out0;
wire v_G2_6350_out0;
wire v_G2_6351_out0;
wire v_G2_6352_out0;
wire v_G2_6353_out0;
wire v_G2_6354_out0;
wire v_G2_6355_out0;
wire v_G2_6356_out0;
wire v_G2_6357_out0;
wire v_G2_6358_out0;
wire v_G2_6359_out0;
wire v_G2_6360_out0;
wire v_G2_6361_out0;
wire v_G2_6362_out0;
wire v_G2_6363_out0;
wire v_G2_6364_out0;
wire v_G2_6365_out0;
wire v_G2_6366_out0;
wire v_G2_6367_out0;
wire v_G2_6368_out0;
wire v_G2_6369_out0;
wire v_G2_6370_out0;
wire v_G2_6371_out0;
wire v_G2_6372_out0;
wire v_G2_6373_out0;
wire v_G2_6374_out0;
wire v_G2_6375_out0;
wire v_G2_6376_out0;
wire v_G2_6377_out0;
wire v_G2_6378_out0;
wire v_G2_6379_out0;
wire v_G2_6380_out0;
wire v_G2_6381_out0;
wire v_G2_6382_out0;
wire v_G2_6383_out0;
wire v_G2_6384_out0;
wire v_G2_6385_out0;
wire v_G2_6386_out0;
wire v_G2_6387_out0;
wire v_G2_6388_out0;
wire v_G2_6389_out0;
wire v_G2_6390_out0;
wire v_G2_6391_out0;
wire v_G2_6392_out0;
wire v_G2_6393_out0;
wire v_G2_6394_out0;
wire v_G2_6395_out0;
wire v_G2_6396_out0;
wire v_G2_6397_out0;
wire v_G2_6398_out0;
wire v_G2_6399_out0;
wire v_G2_6400_out0;
wire v_G2_6401_out0;
wire v_G2_6402_out0;
wire v_G2_6403_out0;
wire v_G2_6404_out0;
wire v_G2_6405_out0;
wire v_G2_6406_out0;
wire v_G2_6407_out0;
wire v_G2_6408_out0;
wire v_G2_6409_out0;
wire v_G2_6410_out0;
wire v_G2_6411_out0;
wire v_G2_6412_out0;
wire v_G2_6413_out0;
wire v_G2_6414_out0;
wire v_G2_6415_out0;
wire v_G2_6416_out0;
wire v_G2_6417_out0;
wire v_G2_6418_out0;
wire v_G2_6419_out0;
wire v_G2_6420_out0;
wire v_G2_6421_out0;
wire v_G2_6422_out0;
wire v_G2_6423_out0;
wire v_G2_6424_out0;
wire v_G2_6425_out0;
wire v_G2_6426_out0;
wire v_G2_6427_out0;
wire v_G2_6428_out0;
wire v_G2_6429_out0;
wire v_G2_6430_out0;
wire v_G2_6431_out0;
wire v_G2_6432_out0;
wire v_G2_6433_out0;
wire v_G2_6434_out0;
wire v_G2_6435_out0;
wire v_G2_6436_out0;
wire v_G2_6437_out0;
wire v_G2_6438_out0;
wire v_G2_6439_out0;
wire v_G2_6440_out0;
wire v_G2_6441_out0;
wire v_G2_6442_out0;
wire v_G2_6443_out0;
wire v_G2_6444_out0;
wire v_G2_6445_out0;
wire v_G2_6446_out0;
wire v_G2_6447_out0;
wire v_G2_6448_out0;
wire v_G2_6449_out0;
wire v_G2_6450_out0;
wire v_G2_6451_out0;
wire v_G2_6452_out0;
wire v_G2_6453_out0;
wire v_G2_6454_out0;
wire v_G2_6455_out0;
wire v_G2_6456_out0;
wire v_G2_6457_out0;
wire v_G2_6458_out0;
wire v_G2_6459_out0;
wire v_G2_6460_out0;
wire v_G2_6461_out0;
wire v_G2_6462_out0;
wire v_G2_6463_out0;
wire v_G2_6464_out0;
wire v_G2_6465_out0;
wire v_G2_6466_out0;
wire v_G2_6467_out0;
wire v_G2_6468_out0;
wire v_G2_6469_out0;
wire v_G2_6470_out0;
wire v_G2_6471_out0;
wire v_G2_6472_out0;
wire v_G2_6473_out0;
wire v_G2_6474_out0;
wire v_G2_6475_out0;
wire v_G2_6476_out0;
wire v_G2_6477_out0;
wire v_G2_6478_out0;
wire v_G2_6479_out0;
wire v_G2_6480_out0;
wire v_G2_6481_out0;
wire v_G2_6482_out0;
wire v_G2_6483_out0;
wire v_G2_6484_out0;
wire v_G2_6485_out0;
wire v_G2_6486_out0;
wire v_G2_6487_out0;
wire v_G2_6488_out0;
wire v_G2_6489_out0;
wire v_G2_6490_out0;
wire v_G2_6491_out0;
wire v_G2_6492_out0;
wire v_G2_6493_out0;
wire v_G2_6494_out0;
wire v_G2_6495_out0;
wire v_G2_6496_out0;
wire v_G2_6497_out0;
wire v_G2_6498_out0;
wire v_G2_6499_out0;
wire v_G2_6723_out0;
wire v_G2_884_out0;
wire v_G2_885_out0;
wire v_G2_923_out0;
wire v_G35_5104_out0;
wire v_G35_5105_out0;
wire v_G36_1528_out0;
wire v_G36_1529_out0;
wire v_G37_3388_out0;
wire v_G37_3389_out0;
wire v_G38_1903_out0;
wire v_G38_1904_out0;
wire v_G3_103_out0;
wire v_G3_104_out0;
wire v_G3_10_out0;
wire v_G3_120_out0;
wire v_G3_121_out0;
wire v_G3_122_out0;
wire v_G3_123_out0;
wire v_G3_124_out0;
wire v_G3_125_out0;
wire v_G3_126_out0;
wire v_G3_1277_out0;
wire v_G3_127_out0;
wire v_G3_128_out0;
wire v_G3_129_out0;
wire v_G3_130_out0;
wire v_G3_1313_out0;
wire v_G3_131_out0;
wire v_G3_132_out0;
wire v_G3_133_out0;
wire v_G3_134_out0;
wire v_G3_1414_out0;
wire v_G3_1435_out0;
wire v_G3_1625_out0;
wire v_G3_1858_out0;
wire v_G3_1932_out0;
wire v_G3_3385_out0;
wire v_G3_3386_out0;
wire v_G3_3479_out0;
wire v_G3_3480_out0;
wire v_G3_4265_out0;
wire v_G3_5151_out0;
wire v_G3_5370_out0;
wire v_G3_6656_out0;
wire v_G3_6720_out0;
wire v_G3_843_out0;
wire v_G3_953_out0;
wire v_G4_109_out0;
wire v_G4_1350_out0;
wire v_G4_1351_out0;
wire v_G4_1575_out0;
wire v_G4_169_out0;
wire v_G4_170_out0;
wire v_G4_171_out0;
wire v_G4_172_out0;
wire v_G4_173_out0;
wire v_G4_174_out0;
wire v_G4_175_out0;
wire v_G4_176_out0;
wire v_G4_177_out0;
wire v_G4_178_out0;
wire v_G4_179_out0;
wire v_G4_180_out0;
wire v_G4_181_out0;
wire v_G4_182_out0;
wire v_G4_183_out0;
wire v_G4_2313_out0;
wire v_G4_2365_out0;
wire v_G4_3394_out0;
wire v_G4_5071_out0;
wire v_G4_5412_out0;
wire v_G4_5413_out0;
wire v_G4_6030_out0;
wire v_G4_6032_out0;
wire v_G4_6750_out0;
wire v_G4_958_out0;
wire v_G4_959_out0;
wire v_G5_102_out0;
wire v_G5_114_out0;
wire v_G5_1260_out0;
wire v_G5_1261_out0;
wire v_G5_1358_out0;
wire v_G5_1359_out0;
wire v_G5_2187_out0;
wire v_G5_221_out0;
wire v_G5_2253_out0;
wire v_G5_309_out0;
wire v_G5_3486_out0;
wire v_G5_5142_out0;
wire v_G5_5183_out0;
wire v_G5_5200_out0;
wire v_G5_5201_out0;
wire v_G5_5228_out0;
wire v_G5_5229_out0;
wire v_G5_5230_out0;
wire v_G5_5231_out0;
wire v_G5_5232_out0;
wire v_G5_5233_out0;
wire v_G5_5234_out0;
wire v_G5_5235_out0;
wire v_G5_5236_out0;
wire v_G5_5237_out0;
wire v_G5_5238_out0;
wire v_G5_5239_out0;
wire v_G5_5240_out0;
wire v_G5_5241_out0;
wire v_G5_5242_out0;
wire v_G5_5369_out0;
wire v_G5_5408_out0;
wire v_G5_587_out0;
wire v_G6_1030_out0;
wire v_G6_1031_out0;
wire v_G6_1032_out0;
wire v_G6_1033_out0;
wire v_G6_1034_out0;
wire v_G6_1035_out0;
wire v_G6_1036_out0;
wire v_G6_1037_out0;
wire v_G6_1038_out0;
wire v_G6_1039_out0;
wire v_G6_1040_out0;
wire v_G6_1041_out0;
wire v_G6_1042_out0;
wire v_G6_1043_out0;
wire v_G6_1044_out0;
wire v_G6_1178_out0;
wire v_G6_1415_out0;
wire v_G6_162_out0;
wire v_G6_2214_out0;
wire v_G6_3443_out0;
wire v_G6_4346_out0;
wire v_G6_4347_out0;
wire v_G6_5508_out0;
wire v_G6_569_out0;
wire v_G6_570_out0;
wire v_G6_6537_out0;
wire v_G6_6648_out0;
wire v_G6_6718_out0;
wire v_G6_6719_out0;
wire v_G7_1195_out0;
wire v_G7_1356_out0;
wire v_G7_1357_out0;
wire v_G7_17_out0;
wire v_G7_2186_out0;
wire v_G7_2354_out0;
wire v_G7_4260_out0;
wire v_G7_4261_out0;
wire v_G7_5093_out0;
wire v_G7_5543_out0;
wire v_G7_5544_out0;
wire v_G7_5545_out0;
wire v_G7_5546_out0;
wire v_G7_5547_out0;
wire v_G7_5548_out0;
wire v_G7_5549_out0;
wire v_G7_5550_out0;
wire v_G7_5551_out0;
wire v_G7_5552_out0;
wire v_G7_5553_out0;
wire v_G7_5554_out0;
wire v_G7_5555_out0;
wire v_G7_5556_out0;
wire v_G7_5557_out0;
wire v_G7_586_out0;
wire v_G7_826_out0;
wire v_G7_87_out0;
wire v_G8_1205_out0;
wire v_G8_1206_out0;
wire v_G8_1207_out0;
wire v_G8_1208_out0;
wire v_G8_1209_out0;
wire v_G8_1210_out0;
wire v_G8_1211_out0;
wire v_G8_1212_out0;
wire v_G8_1213_out0;
wire v_G8_1214_out0;
wire v_G8_1215_out0;
wire v_G8_1216_out0;
wire v_G8_1217_out0;
wire v_G8_1218_out0;
wire v_G8_1219_out0;
wire v_G8_1278_out0;
wire v_G8_1289_out0;
wire v_G8_2178_out0;
wire v_G8_269_out0;
wire v_G8_270_out0;
wire v_G8_5222_out0;
wire v_G8_5223_out0;
wire v_G8_595_out0;
wire v_G8_596_out0;
wire v_G8_6721_out0;
wire v_G8_863_out0;
wire v_G8_987_out0;
wire v_G8_9_out0;
wire v_G9_1046_out0;
wire v_G9_111_out0;
wire v_G9_1138_out0;
wire v_G9_1410_out0;
wire v_G9_1411_out0;
wire v_G9_197_out0;
wire v_G9_199_out0;
wire v_G9_5075_out0;
wire v_G9_5076_out0;
wire v_G9_5203_out0;
wire v_G9_5204_out0;
wire v_G9_5205_out0;
wire v_G9_5206_out0;
wire v_G9_5207_out0;
wire v_G9_5208_out0;
wire v_G9_5209_out0;
wire v_G9_5210_out0;
wire v_G9_5211_out0;
wire v_G9_5212_out0;
wire v_G9_5213_out0;
wire v_G9_5214_out0;
wire v_G9_5215_out0;
wire v_G9_5216_out0;
wire v_G9_5217_out0;
wire v_G9_6551_out0;
wire v_G9_6552_out0;
wire v_G9_6684_out0;
wire v_G9_821_out0;
wire v_INSTRUCTION_32_out0;
wire v_IN_1202_out0;
wire v_IR15_1201_out0;
wire v_JEQZ_1455_out0;
wire v_JEQZ_5174_out0;
wire v_JEQ_1089_out0;
wire v_JEQ_2174_out0;
wire v_JEQ_4334_out0;
wire v_JEQ_5167_out0;
wire v_JEQ_6682_out0;
wire v_JMIN_1298_out0;
wire v_JMIN_590_out0;
wire v_JMI_1565_out0;
wire v_JMI_4273_out0;
wire v_JMI_47_out0;
wire v_JMI_6575_out0;
wire v_JMI_948_out0;
wire v_JMP_1301_out0;
wire v_JMP_1574_out0;
wire v_JMP_268_out0;
wire v_JMP_3475_out0;
wire v_JMP_4342_out0;
wire v_JUMP_1066_out0;
wire v_LOAD_115_out0;
wire v_LOAD_1412_out0;
wire v_LOAD_1519_out0;
wire v_LOAD_3488_out0;
wire v_LOAD_4312_out0;
wire v_LSL_1388_out0;
wire v_LSL_1486_out0;
wire v_LSL_1551_out0;
wire v_LSL_909_out0;
wire v_LSR_204_out0;
wire v_LSR_3393_out0;
wire v_LSR_576_out0;
wire v_LSR_6568_out0;
wire v_MI_1273_out0;
wire v_MI_274_out0;
wire v_MI_5330_out0;
wire v_MOV_5117_out0;
wire v_MOV_99_out0;
wire v_MULTI_INSTRUCTION_1193_out0;
wire v_MULTI_INSTRUCTION_1928_out0;
wire v_MULTI_INSTRUCTION_300_out0;
wire v_MULTI_INSTRUCTION_6558_out0;
wire v_MULTI_INSTRUCTION_6565_out0;
wire v_MULTI_OPCODE_1474_out0;
wire v_MULTI_OPCODE_5461_out0;
wire v_MUX1_1279_out0;
wire v_MUX1_314_out0;
wire v_MUX2_2175_out0;
wire v_MUX3_3503_out0;
wire v_MUX3_4339_out0;
wire v_MUX4_1568_out0;
wire v_MUX5_5060_out0;
wire v_MUX5_6574_out0;
wire v_MUX6_4309_out0;
wire v_MUX6_5401_out0;
wire v_MUX7_5145_out0;
wire v_MUX8_1316_out0;
wire v_MUX9_85_out0;
wire v_NEGATIVE_5541_out0;
wire v_NORMAL_5057_out0;
wire v_NORMAL_6615_out0;
wire v_NORMAL_93_out0;
wire v_NOTUSED1_5259_out0;
wire v_NOTUSED2_2839_out0;
wire v_NOTUSED3_5192_out0;
wire v_NOTUSED4_5182_out0;
wire v_NOTUSED_161_out0;
wire v_NOTUSED_2183_out0;
wire v_NOTUSED_2250_out0;
wire v_NOTUSED_5331_out0;
wire v_NOTUSED_962_out0;
wire v_OP2_SIGN_5333_out0;
wire v_OP2_SIGN_5516_out0;
wire v_OUTSTREAM_1024_out0;
wire v_OUT_13_out0;
wire v_OVERFLOW_5165_out0;
wire v_OVERFLOW_RX_858_out0;
wire v_P_5258_out0;
wire v_Q0_2184_out0;
wire v_Q0_2185_out0;
wire v_Q0_303_out0;
wire v_Q0_5512_out0;
wire v_Q0_5513_out0;
wire v_Q0_6576_out0;
wire v_Q1_1028_out0;
wire v_Q1_152_out0;
wire v_Q1_3390_out0;
wire v_Q1_3391_out0;
wire v_Q1_4358_out0;
wire v_Q1_4359_out0;
wire v_Q2_3378_out0;
wire v_Q2_3379_out0;
wire v_Q2_823_out0;
wire v_Q2_824_out0;
wire v_Q3_4301_out0;
wire v_Q3_4302_out0;
wire v_Q3_5177_out0;
wire v_Q3_5178_out0;
wire v_Q6_924_out0;
wire v_Q6_925_out0;
wire v_Q7_3382_out0;
wire v_Q7_3383_out0;
wire v_Q_144_out0;
wire v_Q_145_out0;
wire v_Q_146_out0;
wire v_Q_147_out0;
wire v_Q_148_out0;
wire v_Q_149_out0;
wire v_Q_150_out0;
wire v_Q_151_out0;
wire v_Q_3786_out0;
wire v_RAMWEN_5267_out0;
wire v_RDN_1628_out0;
wire v_RDN_2196_out0;
wire v_RDN_2197_out0;
wire v_RDN_2198_out0;
wire v_RDN_2199_out0;
wire v_RDN_2200_out0;
wire v_RDN_2201_out0;
wire v_RDN_2202_out0;
wire v_RDN_2203_out0;
wire v_RDN_2204_out0;
wire v_RDN_2205_out0;
wire v_RDN_2206_out0;
wire v_RDN_2207_out0;
wire v_RDN_2208_out0;
wire v_RDN_2209_out0;
wire v_RDN_2210_out0;
wire v_RD_2872_out0;
wire v_RD_2873_out0;
wire v_RD_2874_out0;
wire v_RD_2875_out0;
wire v_RD_2876_out0;
wire v_RD_2877_out0;
wire v_RD_2878_out0;
wire v_RD_2879_out0;
wire v_RD_2880_out0;
wire v_RD_2881_out0;
wire v_RD_2882_out0;
wire v_RD_2883_out0;
wire v_RD_2884_out0;
wire v_RD_2885_out0;
wire v_RD_2886_out0;
wire v_RD_2887_out0;
wire v_RD_2888_out0;
wire v_RD_2889_out0;
wire v_RD_2890_out0;
wire v_RD_2891_out0;
wire v_RD_2892_out0;
wire v_RD_2893_out0;
wire v_RD_2894_out0;
wire v_RD_2895_out0;
wire v_RD_2896_out0;
wire v_RD_2897_out0;
wire v_RD_2898_out0;
wire v_RD_2899_out0;
wire v_RD_2900_out0;
wire v_RD_2901_out0;
wire v_RD_2902_out0;
wire v_RD_2903_out0;
wire v_RD_2904_out0;
wire v_RD_2905_out0;
wire v_RD_2906_out0;
wire v_RD_2907_out0;
wire v_RD_2908_out0;
wire v_RD_2909_out0;
wire v_RD_2910_out0;
wire v_RD_2911_out0;
wire v_RD_2912_out0;
wire v_RD_2913_out0;
wire v_RD_2914_out0;
wire v_RD_2915_out0;
wire v_RD_2916_out0;
wire v_RD_2917_out0;
wire v_RD_2918_out0;
wire v_RD_2919_out0;
wire v_RD_2920_out0;
wire v_RD_2921_out0;
wire v_RD_2922_out0;
wire v_RD_2923_out0;
wire v_RD_2924_out0;
wire v_RD_2925_out0;
wire v_RD_2926_out0;
wire v_RD_2927_out0;
wire v_RD_2928_out0;
wire v_RD_2929_out0;
wire v_RD_2930_out0;
wire v_RD_2931_out0;
wire v_RD_2932_out0;
wire v_RD_2933_out0;
wire v_RD_2934_out0;
wire v_RD_2935_out0;
wire v_RD_2936_out0;
wire v_RD_2937_out0;
wire v_RD_2938_out0;
wire v_RD_2939_out0;
wire v_RD_2940_out0;
wire v_RD_2941_out0;
wire v_RD_2942_out0;
wire v_RD_2943_out0;
wire v_RD_2944_out0;
wire v_RD_2945_out0;
wire v_RD_2946_out0;
wire v_RD_2947_out0;
wire v_RD_2948_out0;
wire v_RD_2949_out0;
wire v_RD_2950_out0;
wire v_RD_2951_out0;
wire v_RD_2952_out0;
wire v_RD_2953_out0;
wire v_RD_2954_out0;
wire v_RD_2955_out0;
wire v_RD_2956_out0;
wire v_RD_2957_out0;
wire v_RD_2958_out0;
wire v_RD_2959_out0;
wire v_RD_2960_out0;
wire v_RD_2961_out0;
wire v_RD_2962_out0;
wire v_RD_2963_out0;
wire v_RD_2964_out0;
wire v_RD_2965_out0;
wire v_RD_2966_out0;
wire v_RD_2967_out0;
wire v_RD_2968_out0;
wire v_RD_2969_out0;
wire v_RD_2970_out0;
wire v_RD_2971_out0;
wire v_RD_2972_out0;
wire v_RD_2973_out0;
wire v_RD_2974_out0;
wire v_RD_2975_out0;
wire v_RD_2976_out0;
wire v_RD_2977_out0;
wire v_RD_2978_out0;
wire v_RD_2979_out0;
wire v_RD_2980_out0;
wire v_RD_2981_out0;
wire v_RD_2982_out0;
wire v_RD_2983_out0;
wire v_RD_2984_out0;
wire v_RD_2985_out0;
wire v_RD_2986_out0;
wire v_RD_2987_out0;
wire v_RD_2988_out0;
wire v_RD_2989_out0;
wire v_RD_2990_out0;
wire v_RD_2991_out0;
wire v_RD_2992_out0;
wire v_RD_2993_out0;
wire v_RD_2994_out0;
wire v_RD_2995_out0;
wire v_RD_2996_out0;
wire v_RD_2997_out0;
wire v_RD_2998_out0;
wire v_RD_2999_out0;
wire v_RD_3000_out0;
wire v_RD_3001_out0;
wire v_RD_3002_out0;
wire v_RD_3003_out0;
wire v_RD_3004_out0;
wire v_RD_3005_out0;
wire v_RD_3006_out0;
wire v_RD_3007_out0;
wire v_RD_3008_out0;
wire v_RD_3009_out0;
wire v_RD_3010_out0;
wire v_RD_3011_out0;
wire v_RD_3012_out0;
wire v_RD_3013_out0;
wire v_RD_3014_out0;
wire v_RD_3015_out0;
wire v_RD_3016_out0;
wire v_RD_3017_out0;
wire v_RD_3018_out0;
wire v_RD_3019_out0;
wire v_RD_3020_out0;
wire v_RD_3021_out0;
wire v_RD_3022_out0;
wire v_RD_3023_out0;
wire v_RD_3024_out0;
wire v_RD_3025_out0;
wire v_RD_3026_out0;
wire v_RD_3027_out0;
wire v_RD_3028_out0;
wire v_RD_3029_out0;
wire v_RD_3030_out0;
wire v_RD_3031_out0;
wire v_RD_3032_out0;
wire v_RD_3033_out0;
wire v_RD_3034_out0;
wire v_RD_3035_out0;
wire v_RD_3036_out0;
wire v_RD_3037_out0;
wire v_RD_3038_out0;
wire v_RD_3039_out0;
wire v_RD_3040_out0;
wire v_RD_3041_out0;
wire v_RD_3042_out0;
wire v_RD_3043_out0;
wire v_RD_3044_out0;
wire v_RD_3045_out0;
wire v_RD_3046_out0;
wire v_RD_3047_out0;
wire v_RD_3048_out0;
wire v_RD_3049_out0;
wire v_RD_3050_out0;
wire v_RD_3051_out0;
wire v_RD_3052_out0;
wire v_RD_3053_out0;
wire v_RD_3054_out0;
wire v_RD_3055_out0;
wire v_RD_3056_out0;
wire v_RD_3057_out0;
wire v_RD_3058_out0;
wire v_RD_3059_out0;
wire v_RD_3060_out0;
wire v_RD_3061_out0;
wire v_RD_3062_out0;
wire v_RD_3063_out0;
wire v_RD_3064_out0;
wire v_RD_3065_out0;
wire v_RD_3066_out0;
wire v_RD_3067_out0;
wire v_RD_3068_out0;
wire v_RD_3069_out0;
wire v_RD_3070_out0;
wire v_RD_3071_out0;
wire v_RD_3072_out0;
wire v_RD_3073_out0;
wire v_RD_3074_out0;
wire v_RD_3075_out0;
wire v_RD_3076_out0;
wire v_RD_3077_out0;
wire v_RD_3078_out0;
wire v_RD_3079_out0;
wire v_RD_3080_out0;
wire v_RD_3081_out0;
wire v_RD_3082_out0;
wire v_RD_3083_out0;
wire v_RD_3084_out0;
wire v_RD_3085_out0;
wire v_RD_3086_out0;
wire v_RD_3087_out0;
wire v_RD_3088_out0;
wire v_RD_3089_out0;
wire v_RD_3090_out0;
wire v_RD_3091_out0;
wire v_RD_3092_out0;
wire v_RD_3093_out0;
wire v_RD_3094_out0;
wire v_RD_3095_out0;
wire v_RD_3096_out0;
wire v_RD_3097_out0;
wire v_RD_3098_out0;
wire v_RD_3099_out0;
wire v_RD_3100_out0;
wire v_RD_3101_out0;
wire v_RD_3102_out0;
wire v_RD_3103_out0;
wire v_RD_3104_out0;
wire v_RD_3105_out0;
wire v_RD_3106_out0;
wire v_RD_3107_out0;
wire v_RD_3108_out0;
wire v_RD_3109_out0;
wire v_RD_3110_out0;
wire v_RD_3111_out0;
wire v_RD_3112_out0;
wire v_RD_3113_out0;
wire v_RD_3114_out0;
wire v_RD_3115_out0;
wire v_RD_3116_out0;
wire v_RD_3117_out0;
wire v_RD_3118_out0;
wire v_RD_3119_out0;
wire v_RD_3120_out0;
wire v_RD_3121_out0;
wire v_RD_3122_out0;
wire v_RD_3123_out0;
wire v_RD_3124_out0;
wire v_RD_3125_out0;
wire v_RD_3126_out0;
wire v_RD_3127_out0;
wire v_RD_3128_out0;
wire v_RD_3129_out0;
wire v_RD_3130_out0;
wire v_RD_3131_out0;
wire v_RD_3132_out0;
wire v_RD_3133_out0;
wire v_RD_3134_out0;
wire v_RD_3135_out0;
wire v_RD_3136_out0;
wire v_RD_3137_out0;
wire v_RD_3138_out0;
wire v_RD_3139_out0;
wire v_RD_3140_out0;
wire v_RD_3141_out0;
wire v_RD_3142_out0;
wire v_RD_3143_out0;
wire v_RD_3144_out0;
wire v_RD_3145_out0;
wire v_RD_3146_out0;
wire v_RD_3147_out0;
wire v_RD_3148_out0;
wire v_RD_3149_out0;
wire v_RD_3150_out0;
wire v_RD_3151_out0;
wire v_RD_3152_out0;
wire v_RD_3153_out0;
wire v_RD_3154_out0;
wire v_RD_3155_out0;
wire v_RD_3156_out0;
wire v_RD_3157_out0;
wire v_RD_3158_out0;
wire v_RD_3159_out0;
wire v_RD_3160_out0;
wire v_RD_3161_out0;
wire v_RD_3162_out0;
wire v_RD_3163_out0;
wire v_RD_3164_out0;
wire v_RD_3165_out0;
wire v_RD_3166_out0;
wire v_RD_3167_out0;
wire v_RD_3168_out0;
wire v_RD_3169_out0;
wire v_RD_3170_out0;
wire v_RD_3171_out0;
wire v_RD_3172_out0;
wire v_RD_3173_out0;
wire v_RD_3174_out0;
wire v_RD_3175_out0;
wire v_RD_3176_out0;
wire v_RD_3177_out0;
wire v_RD_3178_out0;
wire v_RD_3179_out0;
wire v_RD_3180_out0;
wire v_RD_3181_out0;
wire v_RD_3182_out0;
wire v_RD_3183_out0;
wire v_RD_3184_out0;
wire v_RD_3185_out0;
wire v_RD_3186_out0;
wire v_RD_3187_out0;
wire v_RD_3188_out0;
wire v_RD_3189_out0;
wire v_RD_3190_out0;
wire v_RD_3191_out0;
wire v_RD_3192_out0;
wire v_RD_3193_out0;
wire v_RD_3194_out0;
wire v_RD_3195_out0;
wire v_RD_3196_out0;
wire v_RD_3197_out0;
wire v_RD_3198_out0;
wire v_RD_3199_out0;
wire v_RD_3200_out0;
wire v_RD_3201_out0;
wire v_RD_3202_out0;
wire v_RD_3203_out0;
wire v_RD_3204_out0;
wire v_RD_3205_out0;
wire v_RD_3206_out0;
wire v_RD_3207_out0;
wire v_RD_3208_out0;
wire v_RD_3209_out0;
wire v_RD_3210_out0;
wire v_RD_3211_out0;
wire v_RD_3212_out0;
wire v_RD_3213_out0;
wire v_RD_3214_out0;
wire v_RD_3215_out0;
wire v_RD_3216_out0;
wire v_RD_3217_out0;
wire v_RD_3218_out0;
wire v_RD_3219_out0;
wire v_RD_3220_out0;
wire v_RD_3221_out0;
wire v_RD_3222_out0;
wire v_RD_3223_out0;
wire v_RD_3224_out0;
wire v_RD_3225_out0;
wire v_RD_3226_out0;
wire v_RD_3227_out0;
wire v_RD_3228_out0;
wire v_RD_3229_out0;
wire v_RD_3230_out0;
wire v_RD_3231_out0;
wire v_RD_3232_out0;
wire v_RD_3233_out0;
wire v_RD_3234_out0;
wire v_RD_3235_out0;
wire v_RD_3236_out0;
wire v_RD_3237_out0;
wire v_RD_3238_out0;
wire v_RD_3239_out0;
wire v_RD_3240_out0;
wire v_RD_3241_out0;
wire v_RD_3242_out0;
wire v_RD_3243_out0;
wire v_RD_3244_out0;
wire v_RD_3245_out0;
wire v_RD_3246_out0;
wire v_RD_3247_out0;
wire v_RD_3248_out0;
wire v_RD_3249_out0;
wire v_RD_3250_out0;
wire v_RD_3251_out0;
wire v_RD_3252_out0;
wire v_RD_3253_out0;
wire v_RD_3254_out0;
wire v_RD_3255_out0;
wire v_RD_3256_out0;
wire v_RD_3257_out0;
wire v_RD_3258_out0;
wire v_RD_3259_out0;
wire v_RD_3260_out0;
wire v_RD_3261_out0;
wire v_RD_3262_out0;
wire v_RD_3263_out0;
wire v_RD_3264_out0;
wire v_RD_3265_out0;
wire v_RD_3266_out0;
wire v_RD_3267_out0;
wire v_RD_3268_out0;
wire v_RD_3269_out0;
wire v_RD_3270_out0;
wire v_RD_3271_out0;
wire v_RD_3272_out0;
wire v_RD_3273_out0;
wire v_RD_3274_out0;
wire v_RD_3275_out0;
wire v_RD_3276_out0;
wire v_RD_3277_out0;
wire v_RD_3278_out0;
wire v_RD_3279_out0;
wire v_RD_3280_out0;
wire v_RD_3281_out0;
wire v_RD_3282_out0;
wire v_RD_3283_out0;
wire v_RD_3284_out0;
wire v_RD_3285_out0;
wire v_RD_3286_out0;
wire v_RD_3287_out0;
wire v_RD_3288_out0;
wire v_RD_3289_out0;
wire v_RD_3290_out0;
wire v_RD_3291_out0;
wire v_RD_3292_out0;
wire v_RD_3293_out0;
wire v_RD_3294_out0;
wire v_RD_3295_out0;
wire v_RD_3296_out0;
wire v_RD_3297_out0;
wire v_RD_3298_out0;
wire v_RD_3299_out0;
wire v_RD_3300_out0;
wire v_RD_3301_out0;
wire v_RD_3302_out0;
wire v_RD_3303_out0;
wire v_RD_3304_out0;
wire v_RD_3305_out0;
wire v_RD_3306_out0;
wire v_RD_3307_out0;
wire v_RD_3308_out0;
wire v_RD_3309_out0;
wire v_RD_3310_out0;
wire v_RD_3311_out0;
wire v_RD_3312_out0;
wire v_RD_3313_out0;
wire v_RD_3314_out0;
wire v_RD_3315_out0;
wire v_RD_3316_out0;
wire v_RD_3317_out0;
wire v_RD_3318_out0;
wire v_RD_3319_out0;
wire v_RD_3320_out0;
wire v_RD_3321_out0;
wire v_RD_3322_out0;
wire v_RD_3323_out0;
wire v_RD_3324_out0;
wire v_RD_3325_out0;
wire v_RD_3326_out0;
wire v_RD_3327_out0;
wire v_RD_3328_out0;
wire v_RD_3329_out0;
wire v_RD_3330_out0;
wire v_RD_3331_out0;
wire v_RD_3332_out0;
wire v_RD_3333_out0;
wire v_RD_3334_out0;
wire v_RD_3335_out0;
wire v_RD_3527_out0;
wire v_RD_3528_out0;
wire v_RD_3529_out0;
wire v_RD_3530_out0;
wire v_RD_3531_out0;
wire v_RD_3532_out0;
wire v_RD_3533_out0;
wire v_RD_3534_out0;
wire v_RD_3535_out0;
wire v_RD_3536_out0;
wire v_RD_3537_out0;
wire v_RD_3538_out0;
wire v_RD_3539_out0;
wire v_RD_3540_out0;
wire v_RD_3541_out0;
wire v_RD_3542_out0;
wire v_RD_3543_out0;
wire v_RD_3544_out0;
wire v_RD_3545_out0;
wire v_RD_3546_out0;
wire v_RD_3547_out0;
wire v_RD_3548_out0;
wire v_RD_3549_out0;
wire v_RD_3550_out0;
wire v_RD_3551_out0;
wire v_RD_3552_out0;
wire v_RD_3553_out0;
wire v_RD_3554_out0;
wire v_RD_3555_out0;
wire v_RD_3556_out0;
wire v_RD_3557_out0;
wire v_RD_3558_out0;
wire v_RD_3559_out0;
wire v_RD_3560_out0;
wire v_RD_3561_out0;
wire v_RD_3562_out0;
wire v_RD_3563_out0;
wire v_RD_3564_out0;
wire v_RD_3565_out0;
wire v_RD_3566_out0;
wire v_RD_3567_out0;
wire v_RD_3568_out0;
wire v_RD_3569_out0;
wire v_RD_3570_out0;
wire v_RD_3571_out0;
wire v_RD_3572_out0;
wire v_RD_3573_out0;
wire v_RD_3574_out0;
wire v_RD_3575_out0;
wire v_RD_3576_out0;
wire v_RD_3577_out0;
wire v_RD_3578_out0;
wire v_RD_3579_out0;
wire v_RD_3580_out0;
wire v_RD_3581_out0;
wire v_RD_3582_out0;
wire v_RD_3583_out0;
wire v_RD_3584_out0;
wire v_RD_3585_out0;
wire v_RD_3586_out0;
wire v_RD_3587_out0;
wire v_RD_3588_out0;
wire v_RD_3589_out0;
wire v_RD_3590_out0;
wire v_RD_3591_out0;
wire v_RD_3592_out0;
wire v_RD_3593_out0;
wire v_RD_3594_out0;
wire v_RD_3595_out0;
wire v_RD_3596_out0;
wire v_RD_3597_out0;
wire v_RD_3598_out0;
wire v_RD_3599_out0;
wire v_RD_3600_out0;
wire v_RD_3601_out0;
wire v_RD_3602_out0;
wire v_RD_3603_out0;
wire v_RD_3604_out0;
wire v_RD_3605_out0;
wire v_RD_3606_out0;
wire v_RD_3607_out0;
wire v_RD_3608_out0;
wire v_RD_3609_out0;
wire v_RD_3610_out0;
wire v_RD_3611_out0;
wire v_RD_3612_out0;
wire v_RD_3613_out0;
wire v_RD_3614_out0;
wire v_RD_3615_out0;
wire v_RD_3616_out0;
wire v_RD_3617_out0;
wire v_RD_3618_out0;
wire v_RD_3619_out0;
wire v_RD_3620_out0;
wire v_RD_3621_out0;
wire v_RD_3622_out0;
wire v_RD_3623_out0;
wire v_RD_3624_out0;
wire v_RD_3625_out0;
wire v_RD_3626_out0;
wire v_RD_3627_out0;
wire v_RD_3628_out0;
wire v_RD_3629_out0;
wire v_RD_3630_out0;
wire v_RD_3631_out0;
wire v_RD_3632_out0;
wire v_RD_3633_out0;
wire v_RD_3634_out0;
wire v_RD_3635_out0;
wire v_RD_3636_out0;
wire v_RD_3637_out0;
wire v_RD_3638_out0;
wire v_RD_3639_out0;
wire v_RD_3640_out0;
wire v_RD_3641_out0;
wire v_RD_3642_out0;
wire v_RD_3643_out0;
wire v_RD_3644_out0;
wire v_RD_3645_out0;
wire v_RD_3646_out0;
wire v_RD_3647_out0;
wire v_RD_3648_out0;
wire v_RD_3649_out0;
wire v_RD_3650_out0;
wire v_RD_3651_out0;
wire v_RD_3652_out0;
wire v_RD_3653_out0;
wire v_RD_3654_out0;
wire v_RD_3655_out0;
wire v_RD_3656_out0;
wire v_RD_3657_out0;
wire v_RD_3658_out0;
wire v_RD_3659_out0;
wire v_RD_3660_out0;
wire v_RD_3661_out0;
wire v_RD_3662_out0;
wire v_RD_3663_out0;
wire v_RD_3664_out0;
wire v_RD_3665_out0;
wire v_RD_3666_out0;
wire v_RD_3667_out0;
wire v_RD_3668_out0;
wire v_RD_3669_out0;
wire v_RD_3670_out0;
wire v_RD_3671_out0;
wire v_RD_3672_out0;
wire v_RD_3673_out0;
wire v_RD_3674_out0;
wire v_RD_3675_out0;
wire v_RD_3676_out0;
wire v_RD_3677_out0;
wire v_RD_3678_out0;
wire v_RD_3679_out0;
wire v_RD_3680_out0;
wire v_RD_3681_out0;
wire v_RD_3682_out0;
wire v_RD_3683_out0;
wire v_RD_3684_out0;
wire v_RD_3685_out0;
wire v_RD_3686_out0;
wire v_RD_3687_out0;
wire v_RD_3688_out0;
wire v_RD_3689_out0;
wire v_RD_3690_out0;
wire v_RD_3691_out0;
wire v_RD_3692_out0;
wire v_RD_3693_out0;
wire v_RD_3694_out0;
wire v_RD_3695_out0;
wire v_RD_3696_out0;
wire v_RD_3697_out0;
wire v_RD_3698_out0;
wire v_RD_3699_out0;
wire v_RD_3700_out0;
wire v_RD_3701_out0;
wire v_RD_3702_out0;
wire v_RD_3703_out0;
wire v_RD_3704_out0;
wire v_RD_3705_out0;
wire v_RD_3706_out0;
wire v_RD_3707_out0;
wire v_RD_3708_out0;
wire v_RD_3709_out0;
wire v_RD_3710_out0;
wire v_RD_3711_out0;
wire v_RD_3712_out0;
wire v_RD_3713_out0;
wire v_RD_3714_out0;
wire v_RD_3715_out0;
wire v_RD_3716_out0;
wire v_RD_3717_out0;
wire v_RD_3718_out0;
wire v_RD_3719_out0;
wire v_RD_3720_out0;
wire v_RD_3721_out0;
wire v_RD_3722_out0;
wire v_RD_3723_out0;
wire v_RD_3724_out0;
wire v_RD_3725_out0;
wire v_RD_3726_out0;
wire v_RD_3727_out0;
wire v_RD_3728_out0;
wire v_RD_3729_out0;
wire v_RD_3730_out0;
wire v_RD_3731_out0;
wire v_RD_3732_out0;
wire v_RD_3733_out0;
wire v_RD_3734_out0;
wire v_RD_3735_out0;
wire v_RD_3736_out0;
wire v_RD_3737_out0;
wire v_RD_3738_out0;
wire v_RD_3739_out0;
wire v_RD_3740_out0;
wire v_RD_3741_out0;
wire v_RD_3742_out0;
wire v_RD_3743_out0;
wire v_RD_3744_out0;
wire v_RD_3745_out0;
wire v_RD_3746_out0;
wire v_RD_3747_out0;
wire v_RD_3748_out0;
wire v_RD_3749_out0;
wire v_RD_3750_out0;
wire v_RD_6686_out0;
wire v_RD_6687_out0;
wire v_RD_6688_out0;
wire v_RD_6689_out0;
wire v_RD_6690_out0;
wire v_RD_6691_out0;
wire v_RD_6692_out0;
wire v_RD_6693_out0;
wire v_RD_6694_out0;
wire v_RD_6695_out0;
wire v_RD_6696_out0;
wire v_RD_6697_out0;
wire v_RD_6698_out0;
wire v_RD_6699_out0;
wire v_RD_6700_out0;
wire v_RD_SIGN_1173_out0;
wire v_RD_SIGN_141_out0;
wire v_RECEIVER_1BIT_42_out0;
wire v_RECEIVING_INSTRUCTION_5497_out0;
wire v_RESET_5499_out0;
wire v_RESET_5500_out0;
wire v_RESET_5501_out0;
wire v_RESET_5502_out0;
wire v_RESET_5503_out0;
wire v_RESET_5504_out0;
wire v_RESET_5505_out0;
wire v_RESET_5506_out0;
wire v_RM_1630_out0;
wire v_RM_1631_out0;
wire v_RM_1632_out0;
wire v_RM_1633_out0;
wire v_RM_1634_out0;
wire v_RM_1635_out0;
wire v_RM_1636_out0;
wire v_RM_1637_out0;
wire v_RM_1638_out0;
wire v_RM_1639_out0;
wire v_RM_1640_out0;
wire v_RM_1641_out0;
wire v_RM_1642_out0;
wire v_RM_1643_out0;
wire v_RM_1644_out0;
wire v_RM_1645_out0;
wire v_RM_1646_out0;
wire v_RM_1647_out0;
wire v_RM_1648_out0;
wire v_RM_1649_out0;
wire v_RM_1650_out0;
wire v_RM_1651_out0;
wire v_RM_1652_out0;
wire v_RM_1653_out0;
wire v_RM_1654_out0;
wire v_RM_1655_out0;
wire v_RM_1656_out0;
wire v_RM_1657_out0;
wire v_RM_1658_out0;
wire v_RM_1659_out0;
wire v_RM_1660_out0;
wire v_RM_1661_out0;
wire v_RM_1662_out0;
wire v_RM_1663_out0;
wire v_RM_1664_out0;
wire v_RM_1665_out0;
wire v_RM_1666_out0;
wire v_RM_1667_out0;
wire v_RM_1668_out0;
wire v_RM_1669_out0;
wire v_RM_1670_out0;
wire v_RM_1671_out0;
wire v_RM_1672_out0;
wire v_RM_1673_out0;
wire v_RM_1674_out0;
wire v_RM_1675_out0;
wire v_RM_1676_out0;
wire v_RM_1677_out0;
wire v_RM_1678_out0;
wire v_RM_1679_out0;
wire v_RM_1680_out0;
wire v_RM_1681_out0;
wire v_RM_1682_out0;
wire v_RM_1683_out0;
wire v_RM_1684_out0;
wire v_RM_1685_out0;
wire v_RM_1686_out0;
wire v_RM_1687_out0;
wire v_RM_1688_out0;
wire v_RM_1689_out0;
wire v_RM_1690_out0;
wire v_RM_1691_out0;
wire v_RM_1692_out0;
wire v_RM_1693_out0;
wire v_RM_1694_out0;
wire v_RM_1695_out0;
wire v_RM_1696_out0;
wire v_RM_1697_out0;
wire v_RM_1698_out0;
wire v_RM_1699_out0;
wire v_RM_1700_out0;
wire v_RM_1701_out0;
wire v_RM_1702_out0;
wire v_RM_1703_out0;
wire v_RM_1704_out0;
wire v_RM_1705_out0;
wire v_RM_1706_out0;
wire v_RM_1707_out0;
wire v_RM_1708_out0;
wire v_RM_1709_out0;
wire v_RM_1710_out0;
wire v_RM_1711_out0;
wire v_RM_1712_out0;
wire v_RM_1713_out0;
wire v_RM_1714_out0;
wire v_RM_1715_out0;
wire v_RM_1716_out0;
wire v_RM_1717_out0;
wire v_RM_1718_out0;
wire v_RM_1719_out0;
wire v_RM_1720_out0;
wire v_RM_1721_out0;
wire v_RM_1722_out0;
wire v_RM_1723_out0;
wire v_RM_1724_out0;
wire v_RM_1725_out0;
wire v_RM_1726_out0;
wire v_RM_1727_out0;
wire v_RM_1728_out0;
wire v_RM_1729_out0;
wire v_RM_1730_out0;
wire v_RM_1731_out0;
wire v_RM_1732_out0;
wire v_RM_1733_out0;
wire v_RM_1734_out0;
wire v_RM_1735_out0;
wire v_RM_1736_out0;
wire v_RM_1737_out0;
wire v_RM_1738_out0;
wire v_RM_1739_out0;
wire v_RM_1740_out0;
wire v_RM_1741_out0;
wire v_RM_1742_out0;
wire v_RM_1743_out0;
wire v_RM_1744_out0;
wire v_RM_1745_out0;
wire v_RM_1746_out0;
wire v_RM_1747_out0;
wire v_RM_1748_out0;
wire v_RM_1749_out0;
wire v_RM_1750_out0;
wire v_RM_1751_out0;
wire v_RM_1752_out0;
wire v_RM_1753_out0;
wire v_RM_1754_out0;
wire v_RM_1755_out0;
wire v_RM_1756_out0;
wire v_RM_1757_out0;
wire v_RM_1758_out0;
wire v_RM_1759_out0;
wire v_RM_1760_out0;
wire v_RM_1761_out0;
wire v_RM_1762_out0;
wire v_RM_1763_out0;
wire v_RM_1764_out0;
wire v_RM_1765_out0;
wire v_RM_1766_out0;
wire v_RM_1767_out0;
wire v_RM_1768_out0;
wire v_RM_1769_out0;
wire v_RM_1770_out0;
wire v_RM_1771_out0;
wire v_RM_1772_out0;
wire v_RM_1773_out0;
wire v_RM_1774_out0;
wire v_RM_1775_out0;
wire v_RM_1776_out0;
wire v_RM_1777_out0;
wire v_RM_1778_out0;
wire v_RM_1779_out0;
wire v_RM_1780_out0;
wire v_RM_1781_out0;
wire v_RM_1782_out0;
wire v_RM_1783_out0;
wire v_RM_1784_out0;
wire v_RM_1785_out0;
wire v_RM_1786_out0;
wire v_RM_1787_out0;
wire v_RM_1788_out0;
wire v_RM_1789_out0;
wire v_RM_1790_out0;
wire v_RM_1791_out0;
wire v_RM_1792_out0;
wire v_RM_1793_out0;
wire v_RM_1794_out0;
wire v_RM_1795_out0;
wire v_RM_1796_out0;
wire v_RM_1797_out0;
wire v_RM_1798_out0;
wire v_RM_1799_out0;
wire v_RM_1800_out0;
wire v_RM_1801_out0;
wire v_RM_1802_out0;
wire v_RM_1803_out0;
wire v_RM_1804_out0;
wire v_RM_1805_out0;
wire v_RM_1806_out0;
wire v_RM_1807_out0;
wire v_RM_1808_out0;
wire v_RM_1809_out0;
wire v_RM_1810_out0;
wire v_RM_1811_out0;
wire v_RM_1812_out0;
wire v_RM_1813_out0;
wire v_RM_1814_out0;
wire v_RM_1815_out0;
wire v_RM_1816_out0;
wire v_RM_1817_out0;
wire v_RM_1818_out0;
wire v_RM_1819_out0;
wire v_RM_1820_out0;
wire v_RM_1821_out0;
wire v_RM_1822_out0;
wire v_RM_1823_out0;
wire v_RM_1824_out0;
wire v_RM_1825_out0;
wire v_RM_1826_out0;
wire v_RM_1827_out0;
wire v_RM_1828_out0;
wire v_RM_1829_out0;
wire v_RM_1830_out0;
wire v_RM_1831_out0;
wire v_RM_1832_out0;
wire v_RM_1833_out0;
wire v_RM_1834_out0;
wire v_RM_1835_out0;
wire v_RM_1836_out0;
wire v_RM_1837_out0;
wire v_RM_1838_out0;
wire v_RM_1839_out0;
wire v_RM_1840_out0;
wire v_RM_1841_out0;
wire v_RM_1842_out0;
wire v_RM_1843_out0;
wire v_RM_1844_out0;
wire v_RM_1845_out0;
wire v_RM_1846_out0;
wire v_RM_1847_out0;
wire v_RM_1848_out0;
wire v_RM_1849_out0;
wire v_RM_1850_out0;
wire v_RM_1851_out0;
wire v_RM_1852_out0;
wire v_RM_1853_out0;
wire v_RM_5563_out0;
wire v_RM_5564_out0;
wire v_RM_5565_out0;
wire v_RM_5566_out0;
wire v_RM_5567_out0;
wire v_RM_5568_out0;
wire v_RM_5569_out0;
wire v_RM_5570_out0;
wire v_RM_5571_out0;
wire v_RM_5572_out0;
wire v_RM_5573_out0;
wire v_RM_5574_out0;
wire v_RM_5575_out0;
wire v_RM_5576_out0;
wire v_RM_5577_out0;
wire v_RM_5578_out0;
wire v_RM_5579_out0;
wire v_RM_5580_out0;
wire v_RM_5581_out0;
wire v_RM_5582_out0;
wire v_RM_5583_out0;
wire v_RM_5584_out0;
wire v_RM_5585_out0;
wire v_RM_5586_out0;
wire v_RM_5587_out0;
wire v_RM_5588_out0;
wire v_RM_5589_out0;
wire v_RM_5590_out0;
wire v_RM_5591_out0;
wire v_RM_5592_out0;
wire v_RM_5593_out0;
wire v_RM_5594_out0;
wire v_RM_5595_out0;
wire v_RM_5596_out0;
wire v_RM_5597_out0;
wire v_RM_5598_out0;
wire v_RM_5599_out0;
wire v_RM_5600_out0;
wire v_RM_5601_out0;
wire v_RM_5602_out0;
wire v_RM_5603_out0;
wire v_RM_5604_out0;
wire v_RM_5605_out0;
wire v_RM_5606_out0;
wire v_RM_5607_out0;
wire v_RM_5608_out0;
wire v_RM_5609_out0;
wire v_RM_5610_out0;
wire v_RM_5611_out0;
wire v_RM_5612_out0;
wire v_RM_5613_out0;
wire v_RM_5614_out0;
wire v_RM_5615_out0;
wire v_RM_5616_out0;
wire v_RM_5617_out0;
wire v_RM_5618_out0;
wire v_RM_5619_out0;
wire v_RM_5620_out0;
wire v_RM_5621_out0;
wire v_RM_5622_out0;
wire v_RM_5623_out0;
wire v_RM_5624_out0;
wire v_RM_5625_out0;
wire v_RM_5626_out0;
wire v_RM_5627_out0;
wire v_RM_5628_out0;
wire v_RM_5629_out0;
wire v_RM_5630_out0;
wire v_RM_5631_out0;
wire v_RM_5632_out0;
wire v_RM_5633_out0;
wire v_RM_5634_out0;
wire v_RM_5635_out0;
wire v_RM_5636_out0;
wire v_RM_5637_out0;
wire v_RM_5638_out0;
wire v_RM_5639_out0;
wire v_RM_5640_out0;
wire v_RM_5641_out0;
wire v_RM_5642_out0;
wire v_RM_5643_out0;
wire v_RM_5644_out0;
wire v_RM_5645_out0;
wire v_RM_5646_out0;
wire v_RM_5647_out0;
wire v_RM_5648_out0;
wire v_RM_5649_out0;
wire v_RM_5650_out0;
wire v_RM_5651_out0;
wire v_RM_5652_out0;
wire v_RM_5653_out0;
wire v_RM_5654_out0;
wire v_RM_5655_out0;
wire v_RM_5656_out0;
wire v_RM_5657_out0;
wire v_RM_5658_out0;
wire v_RM_5659_out0;
wire v_RM_5660_out0;
wire v_RM_5661_out0;
wire v_RM_5662_out0;
wire v_RM_5663_out0;
wire v_RM_5664_out0;
wire v_RM_5665_out0;
wire v_RM_5666_out0;
wire v_RM_5667_out0;
wire v_RM_5668_out0;
wire v_RM_5669_out0;
wire v_RM_5670_out0;
wire v_RM_5671_out0;
wire v_RM_5672_out0;
wire v_RM_5673_out0;
wire v_RM_5674_out0;
wire v_RM_5675_out0;
wire v_RM_5676_out0;
wire v_RM_5677_out0;
wire v_RM_5678_out0;
wire v_RM_5679_out0;
wire v_RM_5680_out0;
wire v_RM_5681_out0;
wire v_RM_5682_out0;
wire v_RM_5683_out0;
wire v_RM_5684_out0;
wire v_RM_5685_out0;
wire v_RM_5686_out0;
wire v_RM_5687_out0;
wire v_RM_5688_out0;
wire v_RM_5689_out0;
wire v_RM_5690_out0;
wire v_RM_5691_out0;
wire v_RM_5692_out0;
wire v_RM_5693_out0;
wire v_RM_5694_out0;
wire v_RM_5695_out0;
wire v_RM_5696_out0;
wire v_RM_5697_out0;
wire v_RM_5698_out0;
wire v_RM_5699_out0;
wire v_RM_5700_out0;
wire v_RM_5701_out0;
wire v_RM_5702_out0;
wire v_RM_5703_out0;
wire v_RM_5704_out0;
wire v_RM_5705_out0;
wire v_RM_5706_out0;
wire v_RM_5707_out0;
wire v_RM_5708_out0;
wire v_RM_5709_out0;
wire v_RM_5710_out0;
wire v_RM_5711_out0;
wire v_RM_5712_out0;
wire v_RM_5713_out0;
wire v_RM_5714_out0;
wire v_RM_5715_out0;
wire v_RM_5716_out0;
wire v_RM_5717_out0;
wire v_RM_5718_out0;
wire v_RM_5719_out0;
wire v_RM_5720_out0;
wire v_RM_5721_out0;
wire v_RM_5722_out0;
wire v_RM_5723_out0;
wire v_RM_5724_out0;
wire v_RM_5725_out0;
wire v_RM_5726_out0;
wire v_RM_5727_out0;
wire v_RM_5728_out0;
wire v_RM_5729_out0;
wire v_RM_5730_out0;
wire v_RM_5731_out0;
wire v_RM_5732_out0;
wire v_RM_5733_out0;
wire v_RM_5734_out0;
wire v_RM_5735_out0;
wire v_RM_5736_out0;
wire v_RM_5737_out0;
wire v_RM_5738_out0;
wire v_RM_5739_out0;
wire v_RM_5740_out0;
wire v_RM_5741_out0;
wire v_RM_5742_out0;
wire v_RM_5743_out0;
wire v_RM_5744_out0;
wire v_RM_5745_out0;
wire v_RM_5746_out0;
wire v_RM_5747_out0;
wire v_RM_5748_out0;
wire v_RM_5749_out0;
wire v_RM_5750_out0;
wire v_RM_5751_out0;
wire v_RM_5752_out0;
wire v_RM_5753_out0;
wire v_RM_5754_out0;
wire v_RM_5755_out0;
wire v_RM_5756_out0;
wire v_RM_5757_out0;
wire v_RM_5758_out0;
wire v_RM_5759_out0;
wire v_RM_5760_out0;
wire v_RM_5761_out0;
wire v_RM_5762_out0;
wire v_RM_5763_out0;
wire v_RM_5764_out0;
wire v_RM_5765_out0;
wire v_RM_5766_out0;
wire v_RM_5767_out0;
wire v_RM_5768_out0;
wire v_RM_5769_out0;
wire v_RM_5770_out0;
wire v_RM_5771_out0;
wire v_RM_5772_out0;
wire v_RM_5773_out0;
wire v_RM_5774_out0;
wire v_RM_5775_out0;
wire v_RM_5776_out0;
wire v_RM_5777_out0;
wire v_RM_5778_out0;
wire v_RM_5779_out0;
wire v_RM_5780_out0;
wire v_RM_5781_out0;
wire v_RM_5782_out0;
wire v_RM_5783_out0;
wire v_RM_5784_out0;
wire v_RM_5785_out0;
wire v_RM_5786_out0;
wire v_RM_5787_out0;
wire v_RM_5788_out0;
wire v_RM_5789_out0;
wire v_RM_5790_out0;
wire v_RM_5791_out0;
wire v_RM_5792_out0;
wire v_RM_5793_out0;
wire v_RM_5794_out0;
wire v_RM_5795_out0;
wire v_RM_5796_out0;
wire v_RM_5797_out0;
wire v_RM_5798_out0;
wire v_RM_5799_out0;
wire v_RM_5800_out0;
wire v_RM_5801_out0;
wire v_RM_5802_out0;
wire v_RM_5803_out0;
wire v_RM_5804_out0;
wire v_RM_5805_out0;
wire v_RM_5806_out0;
wire v_RM_5807_out0;
wire v_RM_5808_out0;
wire v_RM_5809_out0;
wire v_RM_5810_out0;
wire v_RM_5811_out0;
wire v_RM_5812_out0;
wire v_RM_5813_out0;
wire v_RM_5814_out0;
wire v_RM_5815_out0;
wire v_RM_5816_out0;
wire v_RM_5817_out0;
wire v_RM_5818_out0;
wire v_RM_5819_out0;
wire v_RM_5820_out0;
wire v_RM_5821_out0;
wire v_RM_5822_out0;
wire v_RM_5823_out0;
wire v_RM_5824_out0;
wire v_RM_5825_out0;
wire v_RM_5826_out0;
wire v_RM_5827_out0;
wire v_RM_5828_out0;
wire v_RM_5829_out0;
wire v_RM_5830_out0;
wire v_RM_5831_out0;
wire v_RM_5832_out0;
wire v_RM_5833_out0;
wire v_RM_5834_out0;
wire v_RM_5835_out0;
wire v_RM_5836_out0;
wire v_RM_5837_out0;
wire v_RM_5838_out0;
wire v_RM_5839_out0;
wire v_RM_5840_out0;
wire v_RM_5841_out0;
wire v_RM_5842_out0;
wire v_RM_5843_out0;
wire v_RM_5844_out0;
wire v_RM_5845_out0;
wire v_RM_5846_out0;
wire v_RM_5847_out0;
wire v_RM_5848_out0;
wire v_RM_5849_out0;
wire v_RM_5850_out0;
wire v_RM_5851_out0;
wire v_RM_5852_out0;
wire v_RM_5853_out0;
wire v_RM_5854_out0;
wire v_RM_5855_out0;
wire v_RM_5856_out0;
wire v_RM_5857_out0;
wire v_RM_5858_out0;
wire v_RM_5859_out0;
wire v_RM_5860_out0;
wire v_RM_5861_out0;
wire v_RM_5862_out0;
wire v_RM_5863_out0;
wire v_RM_5864_out0;
wire v_RM_5865_out0;
wire v_RM_5866_out0;
wire v_RM_5867_out0;
wire v_RM_5868_out0;
wire v_RM_5869_out0;
wire v_RM_5870_out0;
wire v_RM_5871_out0;
wire v_RM_5872_out0;
wire v_RM_5873_out0;
wire v_RM_5874_out0;
wire v_RM_5875_out0;
wire v_RM_5876_out0;
wire v_RM_5877_out0;
wire v_RM_5878_out0;
wire v_RM_5879_out0;
wire v_RM_5880_out0;
wire v_RM_5881_out0;
wire v_RM_5882_out0;
wire v_RM_5883_out0;
wire v_RM_5884_out0;
wire v_RM_5885_out0;
wire v_RM_5886_out0;
wire v_RM_5887_out0;
wire v_RM_5888_out0;
wire v_RM_5889_out0;
wire v_RM_5890_out0;
wire v_RM_5891_out0;
wire v_RM_5892_out0;
wire v_RM_5893_out0;
wire v_RM_5894_out0;
wire v_RM_5895_out0;
wire v_RM_5896_out0;
wire v_RM_5897_out0;
wire v_RM_5898_out0;
wire v_RM_5899_out0;
wire v_RM_5900_out0;
wire v_RM_5901_out0;
wire v_RM_5902_out0;
wire v_RM_5903_out0;
wire v_RM_5904_out0;
wire v_RM_5905_out0;
wire v_RM_5906_out0;
wire v_RM_5907_out0;
wire v_RM_5908_out0;
wire v_RM_5909_out0;
wire v_RM_5910_out0;
wire v_RM_5911_out0;
wire v_RM_5912_out0;
wire v_RM_5913_out0;
wire v_RM_5914_out0;
wire v_RM_5915_out0;
wire v_RM_5916_out0;
wire v_RM_5917_out0;
wire v_RM_5918_out0;
wire v_RM_5919_out0;
wire v_RM_5920_out0;
wire v_RM_5921_out0;
wire v_RM_5922_out0;
wire v_RM_5923_out0;
wire v_RM_5924_out0;
wire v_RM_5925_out0;
wire v_RM_5926_out0;
wire v_RM_5927_out0;
wire v_RM_5928_out0;
wire v_RM_5929_out0;
wire v_RM_5930_out0;
wire v_RM_5931_out0;
wire v_RM_5932_out0;
wire v_RM_5933_out0;
wire v_RM_5934_out0;
wire v_RM_5935_out0;
wire v_RM_5936_out0;
wire v_RM_5937_out0;
wire v_RM_5938_out0;
wire v_RM_5939_out0;
wire v_RM_5940_out0;
wire v_RM_5941_out0;
wire v_RM_5942_out0;
wire v_RM_5943_out0;
wire v_RM_5944_out0;
wire v_RM_5945_out0;
wire v_RM_5946_out0;
wire v_RM_5947_out0;
wire v_RM_5948_out0;
wire v_RM_5949_out0;
wire v_RM_5950_out0;
wire v_RM_5951_out0;
wire v_RM_5952_out0;
wire v_RM_5953_out0;
wire v_RM_5954_out0;
wire v_RM_5955_out0;
wire v_RM_5956_out0;
wire v_RM_5957_out0;
wire v_RM_5958_out0;
wire v_RM_5959_out0;
wire v_RM_5960_out0;
wire v_RM_5961_out0;
wire v_RM_5962_out0;
wire v_RM_5963_out0;
wire v_RM_5964_out0;
wire v_RM_5965_out0;
wire v_RM_5966_out0;
wire v_RM_5967_out0;
wire v_RM_5968_out0;
wire v_RM_5969_out0;
wire v_RM_5970_out0;
wire v_RM_5971_out0;
wire v_RM_5972_out0;
wire v_RM_5973_out0;
wire v_RM_5974_out0;
wire v_RM_5975_out0;
wire v_RM_5976_out0;
wire v_RM_5977_out0;
wire v_RM_5978_out0;
wire v_RM_5979_out0;
wire v_RM_5980_out0;
wire v_RM_5981_out0;
wire v_RM_5982_out0;
wire v_RM_5983_out0;
wire v_RM_5984_out0;
wire v_RM_5985_out0;
wire v_RM_5986_out0;
wire v_RM_5987_out0;
wire v_RM_5988_out0;
wire v_RM_5989_out0;
wire v_RM_5990_out0;
wire v_RM_5991_out0;
wire v_RM_5992_out0;
wire v_RM_5993_out0;
wire v_RM_5994_out0;
wire v_RM_5995_out0;
wire v_RM_5996_out0;
wire v_RM_5997_out0;
wire v_RM_5998_out0;
wire v_RM_5999_out0;
wire v_RM_6000_out0;
wire v_RM_6001_out0;
wire v_RM_6002_out0;
wire v_RM_6003_out0;
wire v_RM_6004_out0;
wire v_RM_6005_out0;
wire v_RM_6006_out0;
wire v_RM_6007_out0;
wire v_RM_6008_out0;
wire v_RM_6009_out0;
wire v_RM_6010_out0;
wire v_RM_6011_out0;
wire v_RM_6012_out0;
wire v_RM_6013_out0;
wire v_RM_6014_out0;
wire v_RM_6015_out0;
wire v_RM_6016_out0;
wire v_RM_6017_out0;
wire v_RM_6018_out0;
wire v_RM_6019_out0;
wire v_RM_6020_out0;
wire v_RM_6021_out0;
wire v_RM_6022_out0;
wire v_RM_6023_out0;
wire v_RM_6024_out0;
wire v_RM_6025_out0;
wire v_RM_6026_out0;
wire v_ROM1_225_out0;
wire v_ROR_140_out0;
wire v_ROR_1598_out0;
wire v_ROR_1599_out0;
wire v_ROR_267_out0;
wire v_RX_INSTRUCTION_1586_out0;
wire v_RX_INST_49_out0;
wire v_RX_OVERFLOW_15_out0;
wire v_RX_OVERFLOW_5535_out0;
wire v_SBC_2356_out0;
wire v_SBC_5438_out0;
wire v_SBC_6705_out0;
wire v_SEL1_1125_out0;
wire v_SEL1_1130_out0;
wire v_SEL1_1183_out0;
wire v_SEL1_119_out0;
wire v_SEL1_2371_out0;
wire v_SEL1_5081_out0;
wire v_SEL1_571_out0;
wire v_SEL1_589_out0;
wire v_SEL1_6622_out0;
wire v_SEL2_5089_out0;
wire v_SEL3_1274_out0;
wire v_SEL3_561_out0;
wire v_SEL4_3752_out0;
wire v_SEL5_1487_out0;
wire v_SHIFHT_ENABLE_6652_out0;
wire v_SHIFHT_ENABLE_6653_out0;
wire v_SHIFT_ENABLE_4275_out0;
wire v_SHIFT_RD_1240_out0;
wire v_SHIFT_WHICH_OP_2181_out0;
wire v_SHIFT_WHICH_OP_5153_out0;
wire v_SHIFT_WHICH_OP_5274_out0;
wire v_SIGN_ANS_2180_out0;
wire v_SIGN_ANS_4257_out0;
wire v_SIGN_ANS_5080_out0;
wire v_SIGN_ANS_963_out0;
wire v_STALL_208_out0;
wire v_STALL_3392_out0;
wire v_STALL_5070_out0;
wire v_STALL_860_out0;
wire v_STARTBIT_3420_out0;
wire v_STARTBIT_3421_out0;
wire v_START_1476_out0;
wire v_START_191_out0;
wire v_START_6598_out0;
wire v_STORE_110_out0;
wire v_STORE_265_out0;
wire v_STORE_5329_out0;
wire v_STORE_585_out0;
wire v_STORE_6555_out0;
wire v_STP_28_out0;
wire v_STP_5101_out0;
wire v_STP_5154_out0;
wire v_STP_5402_out0;
wire v_STP_5531_out0;
wire v_SUBNORMAL_4335_out0;
wire v_SUB_1315_out0;
wire v_SUB_1417_out0;
wire v_SUB_1442_out0;
wire v_SUB_2255_out0;
wire v_SUB_2256_out0;
wire v_SUB_4264_out0;
wire v_SUB_6033_out0;
wire v_SUB_INSTRUCTION_1361_out0;
wire v_SUB_INSTRUCTION_3478_out0;
wire v_SUB_INSTRUCTION_5510_out0;
wire v_S_2278_out0;
wire v_S_2279_out0;
wire v_S_2280_out0;
wire v_S_2281_out0;
wire v_S_2282_out0;
wire v_S_2283_out0;
wire v_S_2284_out0;
wire v_S_2285_out0;
wire v_S_2286_out0;
wire v_S_2287_out0;
wire v_S_2288_out0;
wire v_S_2289_out0;
wire v_S_2290_out0;
wire v_S_2291_out0;
wire v_S_2292_out0;
wire v_S_4360_out0;
wire v_S_4361_out0;
wire v_S_4362_out0;
wire v_S_4363_out0;
wire v_S_4364_out0;
wire v_S_4365_out0;
wire v_S_4366_out0;
wire v_S_4367_out0;
wire v_S_4368_out0;
wire v_S_4369_out0;
wire v_S_4370_out0;
wire v_S_4371_out0;
wire v_S_4372_out0;
wire v_S_4373_out0;
wire v_S_4374_out0;
wire v_S_4375_out0;
wire v_S_4376_out0;
wire v_S_4377_out0;
wire v_S_4378_out0;
wire v_S_4379_out0;
wire v_S_4380_out0;
wire v_S_4381_out0;
wire v_S_4382_out0;
wire v_S_4383_out0;
wire v_S_4384_out0;
wire v_S_4385_out0;
wire v_S_4386_out0;
wire v_S_4387_out0;
wire v_S_4388_out0;
wire v_S_4389_out0;
wire v_S_4390_out0;
wire v_S_4391_out0;
wire v_S_4392_out0;
wire v_S_4393_out0;
wire v_S_4394_out0;
wire v_S_4395_out0;
wire v_S_4396_out0;
wire v_S_4397_out0;
wire v_S_4398_out0;
wire v_S_4399_out0;
wire v_S_4400_out0;
wire v_S_4401_out0;
wire v_S_4402_out0;
wire v_S_4403_out0;
wire v_S_4404_out0;
wire v_S_4405_out0;
wire v_S_4406_out0;
wire v_S_4407_out0;
wire v_S_4408_out0;
wire v_S_4409_out0;
wire v_S_4410_out0;
wire v_S_4411_out0;
wire v_S_4412_out0;
wire v_S_4413_out0;
wire v_S_4414_out0;
wire v_S_4415_out0;
wire v_S_4416_out0;
wire v_S_4417_out0;
wire v_S_4418_out0;
wire v_S_4419_out0;
wire v_S_4420_out0;
wire v_S_4421_out0;
wire v_S_4422_out0;
wire v_S_4423_out0;
wire v_S_4424_out0;
wire v_S_4425_out0;
wire v_S_4426_out0;
wire v_S_4427_out0;
wire v_S_4428_out0;
wire v_S_4429_out0;
wire v_S_4430_out0;
wire v_S_4431_out0;
wire v_S_4432_out0;
wire v_S_4433_out0;
wire v_S_4434_out0;
wire v_S_4435_out0;
wire v_S_4436_out0;
wire v_S_4437_out0;
wire v_S_4438_out0;
wire v_S_4439_out0;
wire v_S_4440_out0;
wire v_S_4441_out0;
wire v_S_4442_out0;
wire v_S_4443_out0;
wire v_S_4444_out0;
wire v_S_4445_out0;
wire v_S_4446_out0;
wire v_S_4447_out0;
wire v_S_4448_out0;
wire v_S_4449_out0;
wire v_S_4450_out0;
wire v_S_4451_out0;
wire v_S_4452_out0;
wire v_S_4453_out0;
wire v_S_4454_out0;
wire v_S_4455_out0;
wire v_S_4456_out0;
wire v_S_4457_out0;
wire v_S_4458_out0;
wire v_S_4459_out0;
wire v_S_4460_out0;
wire v_S_4461_out0;
wire v_S_4462_out0;
wire v_S_4463_out0;
wire v_S_4464_out0;
wire v_S_4465_out0;
wire v_S_4466_out0;
wire v_S_4467_out0;
wire v_S_4468_out0;
wire v_S_4469_out0;
wire v_S_4470_out0;
wire v_S_4471_out0;
wire v_S_4472_out0;
wire v_S_4473_out0;
wire v_S_4474_out0;
wire v_S_4475_out0;
wire v_S_4476_out0;
wire v_S_4477_out0;
wire v_S_4478_out0;
wire v_S_4479_out0;
wire v_S_4480_out0;
wire v_S_4481_out0;
wire v_S_4482_out0;
wire v_S_4483_out0;
wire v_S_4484_out0;
wire v_S_4485_out0;
wire v_S_4486_out0;
wire v_S_4487_out0;
wire v_S_4488_out0;
wire v_S_4489_out0;
wire v_S_4490_out0;
wire v_S_4491_out0;
wire v_S_4492_out0;
wire v_S_4493_out0;
wire v_S_4494_out0;
wire v_S_4495_out0;
wire v_S_4496_out0;
wire v_S_4497_out0;
wire v_S_4498_out0;
wire v_S_4499_out0;
wire v_S_4500_out0;
wire v_S_4501_out0;
wire v_S_4502_out0;
wire v_S_4503_out0;
wire v_S_4504_out0;
wire v_S_4505_out0;
wire v_S_4506_out0;
wire v_S_4507_out0;
wire v_S_4508_out0;
wire v_S_4509_out0;
wire v_S_4510_out0;
wire v_S_4511_out0;
wire v_S_4512_out0;
wire v_S_4513_out0;
wire v_S_4514_out0;
wire v_S_4515_out0;
wire v_S_4516_out0;
wire v_S_4517_out0;
wire v_S_4518_out0;
wire v_S_4519_out0;
wire v_S_4520_out0;
wire v_S_4521_out0;
wire v_S_4522_out0;
wire v_S_4523_out0;
wire v_S_4524_out0;
wire v_S_4525_out0;
wire v_S_4526_out0;
wire v_S_4527_out0;
wire v_S_4528_out0;
wire v_S_4529_out0;
wire v_S_4530_out0;
wire v_S_4531_out0;
wire v_S_4532_out0;
wire v_S_4533_out0;
wire v_S_4534_out0;
wire v_S_4535_out0;
wire v_S_4536_out0;
wire v_S_4537_out0;
wire v_S_4538_out0;
wire v_S_4539_out0;
wire v_S_4540_out0;
wire v_S_4541_out0;
wire v_S_4542_out0;
wire v_S_4543_out0;
wire v_S_4544_out0;
wire v_S_4545_out0;
wire v_S_4546_out0;
wire v_S_4547_out0;
wire v_S_4548_out0;
wire v_S_4549_out0;
wire v_S_4550_out0;
wire v_S_4551_out0;
wire v_S_4552_out0;
wire v_S_4553_out0;
wire v_S_4554_out0;
wire v_S_4555_out0;
wire v_S_4556_out0;
wire v_S_4557_out0;
wire v_S_4558_out0;
wire v_S_4559_out0;
wire v_S_4560_out0;
wire v_S_4561_out0;
wire v_S_4562_out0;
wire v_S_4563_out0;
wire v_S_4564_out0;
wire v_S_4565_out0;
wire v_S_4566_out0;
wire v_S_4567_out0;
wire v_S_4568_out0;
wire v_S_4569_out0;
wire v_S_4570_out0;
wire v_S_4571_out0;
wire v_S_4572_out0;
wire v_S_4573_out0;
wire v_S_4574_out0;
wire v_S_4575_out0;
wire v_S_4576_out0;
wire v_S_4577_out0;
wire v_S_4578_out0;
wire v_S_4579_out0;
wire v_S_4580_out0;
wire v_S_4581_out0;
wire v_S_4582_out0;
wire v_S_4583_out0;
wire v_S_4584_out0;
wire v_S_4585_out0;
wire v_S_4586_out0;
wire v_S_4587_out0;
wire v_S_4588_out0;
wire v_S_4589_out0;
wire v_S_4590_out0;
wire v_S_4591_out0;
wire v_S_4592_out0;
wire v_S_4593_out0;
wire v_S_4594_out0;
wire v_S_4595_out0;
wire v_S_4596_out0;
wire v_S_4597_out0;
wire v_S_4598_out0;
wire v_S_4599_out0;
wire v_S_4600_out0;
wire v_S_4601_out0;
wire v_S_4602_out0;
wire v_S_4603_out0;
wire v_S_4604_out0;
wire v_S_4605_out0;
wire v_S_4606_out0;
wire v_S_4607_out0;
wire v_S_4608_out0;
wire v_S_4609_out0;
wire v_S_4610_out0;
wire v_S_4611_out0;
wire v_S_4612_out0;
wire v_S_4613_out0;
wire v_S_4614_out0;
wire v_S_4615_out0;
wire v_S_4616_out0;
wire v_S_4617_out0;
wire v_S_4618_out0;
wire v_S_4619_out0;
wire v_S_4620_out0;
wire v_S_4621_out0;
wire v_S_4622_out0;
wire v_S_4623_out0;
wire v_S_4624_out0;
wire v_S_4625_out0;
wire v_S_4626_out0;
wire v_S_4627_out0;
wire v_S_4628_out0;
wire v_S_4629_out0;
wire v_S_4630_out0;
wire v_S_4631_out0;
wire v_S_4632_out0;
wire v_S_4633_out0;
wire v_S_4634_out0;
wire v_S_4635_out0;
wire v_S_4636_out0;
wire v_S_4637_out0;
wire v_S_4638_out0;
wire v_S_4639_out0;
wire v_S_4640_out0;
wire v_S_4641_out0;
wire v_S_4642_out0;
wire v_S_4643_out0;
wire v_S_4644_out0;
wire v_S_4645_out0;
wire v_S_4646_out0;
wire v_S_4647_out0;
wire v_S_4648_out0;
wire v_S_4649_out0;
wire v_S_4650_out0;
wire v_S_4651_out0;
wire v_S_4652_out0;
wire v_S_4653_out0;
wire v_S_4654_out0;
wire v_S_4655_out0;
wire v_S_4656_out0;
wire v_S_4657_out0;
wire v_S_4658_out0;
wire v_S_4659_out0;
wire v_S_4660_out0;
wire v_S_4661_out0;
wire v_S_4662_out0;
wire v_S_4663_out0;
wire v_S_4664_out0;
wire v_S_4665_out0;
wire v_S_4666_out0;
wire v_S_4667_out0;
wire v_S_4668_out0;
wire v_S_4669_out0;
wire v_S_4670_out0;
wire v_S_4671_out0;
wire v_S_4672_out0;
wire v_S_4673_out0;
wire v_S_4674_out0;
wire v_S_4675_out0;
wire v_S_4676_out0;
wire v_S_4677_out0;
wire v_S_4678_out0;
wire v_S_4679_out0;
wire v_S_4680_out0;
wire v_S_4681_out0;
wire v_S_4682_out0;
wire v_S_4683_out0;
wire v_S_4684_out0;
wire v_S_4685_out0;
wire v_S_4686_out0;
wire v_S_4687_out0;
wire v_S_4688_out0;
wire v_S_4689_out0;
wire v_S_4690_out0;
wire v_S_4691_out0;
wire v_S_4692_out0;
wire v_S_4693_out0;
wire v_S_4694_out0;
wire v_S_4695_out0;
wire v_S_4696_out0;
wire v_S_4697_out0;
wire v_S_4698_out0;
wire v_S_4699_out0;
wire v_S_4700_out0;
wire v_S_4701_out0;
wire v_S_4702_out0;
wire v_S_4703_out0;
wire v_S_4704_out0;
wire v_S_4705_out0;
wire v_S_4706_out0;
wire v_S_4707_out0;
wire v_S_4708_out0;
wire v_S_4709_out0;
wire v_S_4710_out0;
wire v_S_4711_out0;
wire v_S_4712_out0;
wire v_S_4713_out0;
wire v_S_4714_out0;
wire v_S_4715_out0;
wire v_S_4716_out0;
wire v_S_4717_out0;
wire v_S_4718_out0;
wire v_S_4719_out0;
wire v_S_4720_out0;
wire v_S_4721_out0;
wire v_S_4722_out0;
wire v_S_4723_out0;
wire v_S_4724_out0;
wire v_S_4725_out0;
wire v_S_4726_out0;
wire v_S_4727_out0;
wire v_S_4728_out0;
wire v_S_4729_out0;
wire v_S_4730_out0;
wire v_S_4731_out0;
wire v_S_4732_out0;
wire v_S_4733_out0;
wire v_S_4734_out0;
wire v_S_4735_out0;
wire v_S_4736_out0;
wire v_S_4737_out0;
wire v_S_4738_out0;
wire v_S_4739_out0;
wire v_S_4740_out0;
wire v_S_4741_out0;
wire v_S_4742_out0;
wire v_S_4743_out0;
wire v_S_4744_out0;
wire v_S_4745_out0;
wire v_S_4746_out0;
wire v_S_4747_out0;
wire v_S_4748_out0;
wire v_S_4749_out0;
wire v_S_4750_out0;
wire v_S_4751_out0;
wire v_S_4752_out0;
wire v_S_4753_out0;
wire v_S_4754_out0;
wire v_S_4755_out0;
wire v_S_4756_out0;
wire v_S_4757_out0;
wire v_S_4758_out0;
wire v_S_4759_out0;
wire v_S_4760_out0;
wire v_S_4761_out0;
wire v_S_4762_out0;
wire v_S_4763_out0;
wire v_S_4764_out0;
wire v_S_4765_out0;
wire v_S_4766_out0;
wire v_S_4767_out0;
wire v_S_4768_out0;
wire v_S_4769_out0;
wire v_S_4770_out0;
wire v_S_4771_out0;
wire v_S_4772_out0;
wire v_S_4773_out0;
wire v_S_4774_out0;
wire v_S_4775_out0;
wire v_S_4776_out0;
wire v_S_4777_out0;
wire v_S_4778_out0;
wire v_S_4779_out0;
wire v_S_4780_out0;
wire v_S_4781_out0;
wire v_S_4782_out0;
wire v_S_4783_out0;
wire v_S_4784_out0;
wire v_S_4785_out0;
wire v_S_4786_out0;
wire v_S_4787_out0;
wire v_S_4788_out0;
wire v_S_4789_out0;
wire v_S_4790_out0;
wire v_S_4791_out0;
wire v_S_4792_out0;
wire v_S_4793_out0;
wire v_S_4794_out0;
wire v_S_4795_out0;
wire v_S_4796_out0;
wire v_S_4797_out0;
wire v_S_4798_out0;
wire v_S_4799_out0;
wire v_S_4800_out0;
wire v_S_4801_out0;
wire v_S_4802_out0;
wire v_S_4803_out0;
wire v_S_4804_out0;
wire v_S_4805_out0;
wire v_S_4806_out0;
wire v_S_4807_out0;
wire v_S_4808_out0;
wire v_S_4809_out0;
wire v_S_4810_out0;
wire v_S_4811_out0;
wire v_S_4812_out0;
wire v_S_4813_out0;
wire v_S_4814_out0;
wire v_S_4815_out0;
wire v_S_4816_out0;
wire v_S_4817_out0;
wire v_S_4818_out0;
wire v_S_4819_out0;
wire v_S_4820_out0;
wire v_S_4821_out0;
wire v_S_4822_out0;
wire v_S_4823_out0;
wire v_S_5562_out0;
wire v_S_597_out0;
wire v_S_598_out0;
wire v_S_599_out0;
wire v_S_600_out0;
wire v_S_601_out0;
wire v_S_602_out0;
wire v_S_603_out0;
wire v_S_604_out0;
wire v_S_605_out0;
wire v_S_606_out0;
wire v_S_607_out0;
wire v_S_608_out0;
wire v_S_609_out0;
wire v_S_610_out0;
wire v_S_611_out0;
wire v_S_612_out0;
wire v_S_613_out0;
wire v_S_614_out0;
wire v_S_615_out0;
wire v_S_616_out0;
wire v_S_617_out0;
wire v_S_618_out0;
wire v_S_619_out0;
wire v_S_620_out0;
wire v_S_621_out0;
wire v_S_622_out0;
wire v_S_623_out0;
wire v_S_624_out0;
wire v_S_625_out0;
wire v_S_626_out0;
wire v_S_627_out0;
wire v_S_628_out0;
wire v_S_629_out0;
wire v_S_630_out0;
wire v_S_631_out0;
wire v_S_632_out0;
wire v_S_633_out0;
wire v_S_634_out0;
wire v_S_635_out0;
wire v_S_636_out0;
wire v_S_637_out0;
wire v_S_638_out0;
wire v_S_639_out0;
wire v_S_640_out0;
wire v_S_641_out0;
wire v_S_642_out0;
wire v_S_643_out0;
wire v_S_644_out0;
wire v_S_645_out0;
wire v_S_646_out0;
wire v_S_647_out0;
wire v_S_648_out0;
wire v_S_649_out0;
wire v_S_650_out0;
wire v_S_651_out0;
wire v_S_652_out0;
wire v_S_653_out0;
wire v_S_654_out0;
wire v_S_655_out0;
wire v_S_656_out0;
wire v_S_657_out0;
wire v_S_658_out0;
wire v_S_659_out0;
wire v_S_660_out0;
wire v_S_661_out0;
wire v_S_662_out0;
wire v_S_663_out0;
wire v_S_664_out0;
wire v_S_665_out0;
wire v_S_666_out0;
wire v_S_667_out0;
wire v_S_668_out0;
wire v_S_669_out0;
wire v_S_670_out0;
wire v_S_671_out0;
wire v_S_672_out0;
wire v_S_673_out0;
wire v_S_674_out0;
wire v_S_675_out0;
wire v_S_676_out0;
wire v_S_677_out0;
wire v_S_678_out0;
wire v_S_679_out0;
wire v_S_680_out0;
wire v_S_681_out0;
wire v_S_682_out0;
wire v_S_683_out0;
wire v_S_684_out0;
wire v_S_685_out0;
wire v_S_686_out0;
wire v_S_687_out0;
wire v_S_688_out0;
wire v_S_689_out0;
wire v_S_690_out0;
wire v_S_691_out0;
wire v_S_692_out0;
wire v_S_693_out0;
wire v_S_694_out0;
wire v_S_695_out0;
wire v_S_696_out0;
wire v_S_697_out0;
wire v_S_698_out0;
wire v_S_699_out0;
wire v_S_700_out0;
wire v_S_701_out0;
wire v_S_702_out0;
wire v_S_703_out0;
wire v_S_704_out0;
wire v_S_705_out0;
wire v_S_706_out0;
wire v_S_707_out0;
wire v_S_708_out0;
wire v_S_709_out0;
wire v_S_710_out0;
wire v_S_711_out0;
wire v_S_712_out0;
wire v_S_713_out0;
wire v_S_714_out0;
wire v_S_715_out0;
wire v_S_716_out0;
wire v_S_717_out0;
wire v_S_718_out0;
wire v_S_719_out0;
wire v_S_720_out0;
wire v_S_721_out0;
wire v_S_722_out0;
wire v_S_723_out0;
wire v_S_724_out0;
wire v_S_725_out0;
wire v_S_726_out0;
wire v_S_727_out0;
wire v_S_728_out0;
wire v_S_729_out0;
wire v_S_730_out0;
wire v_S_731_out0;
wire v_S_732_out0;
wire v_S_733_out0;
wire v_S_734_out0;
wire v_S_735_out0;
wire v_S_736_out0;
wire v_S_737_out0;
wire v_S_738_out0;
wire v_S_739_out0;
wire v_S_740_out0;
wire v_S_741_out0;
wire v_S_742_out0;
wire v_S_743_out0;
wire v_S_744_out0;
wire v_S_745_out0;
wire v_S_746_out0;
wire v_S_747_out0;
wire v_S_748_out0;
wire v_S_749_out0;
wire v_S_750_out0;
wire v_S_751_out0;
wire v_S_752_out0;
wire v_S_753_out0;
wire v_S_754_out0;
wire v_S_755_out0;
wire v_S_756_out0;
wire v_S_757_out0;
wire v_S_758_out0;
wire v_S_759_out0;
wire v_S_760_out0;
wire v_S_761_out0;
wire v_S_762_out0;
wire v_S_763_out0;
wire v_S_764_out0;
wire v_S_765_out0;
wire v_S_766_out0;
wire v_S_767_out0;
wire v_S_768_out0;
wire v_S_769_out0;
wire v_S_770_out0;
wire v_S_771_out0;
wire v_S_772_out0;
wire v_S_773_out0;
wire v_S_774_out0;
wire v_S_775_out0;
wire v_S_776_out0;
wire v_S_777_out0;
wire v_S_778_out0;
wire v_S_779_out0;
wire v_S_780_out0;
wire v_S_781_out0;
wire v_S_782_out0;
wire v_S_783_out0;
wire v_S_784_out0;
wire v_S_785_out0;
wire v_S_786_out0;
wire v_S_787_out0;
wire v_S_788_out0;
wire v_S_789_out0;
wire v_S_790_out0;
wire v_S_791_out0;
wire v_S_792_out0;
wire v_S_793_out0;
wire v_S_794_out0;
wire v_S_795_out0;
wire v_S_796_out0;
wire v_S_797_out0;
wire v_S_798_out0;
wire v_S_799_out0;
wire v_S_800_out0;
wire v_S_801_out0;
wire v_S_802_out0;
wire v_S_803_out0;
wire v_S_804_out0;
wire v_S_805_out0;
wire v_S_806_out0;
wire v_S_807_out0;
wire v_S_808_out0;
wire v_S_809_out0;
wire v_S_810_out0;
wire v_S_811_out0;
wire v_S_812_out0;
wire v_S_813_out0;
wire v_S_814_out0;
wire v_S_815_out0;
wire v_S_816_out0;
wire v_S_817_out0;
wire v_S_818_out0;
wire v_S_819_out0;
wire v_S_820_out0;
wire v_TRANSMITER_1BIT_1200_out0;
wire v_TRANSMITER_OVERFLOW_4268_out0;
wire v_TRANSMITER_OVERFLOW_830_out0;
wire v_TRANSMIT_INSTRUCTION_839_out0;
wire v_TST_1861_out0;
wire v_TST_198_out0;
wire v_TST_4300_out0;
wire v_TX_INSTRUCTION_3442_out0;
wire v_TX_IN_PROGRESS_911_out0;
wire v_TX_IN_PROG_5059_out0;
wire v_TX_OVERFLOW_1902_out0;
wire v_UART_1897_out0;
wire v_UART_5176_out0;
wire v_UART_5325_out0;
wire v_UART_890_out0;
wire v_UNDERFLOW_3395_out0;
wire v_UNNOTUSED_5522_out0;
wire v_UNUSED1_1472_out0;
wire v_UNUSED2_1069_out0;
wire v_UNUSED_168_out0;
wire v_U_5155_out0;
wire v_WEN3_829_out0;
wire v_WENALU_4262_out0;
wire v_WENALU_5345_out0;
wire v_WENLDST_1309_out0;
wire v_WENLDST_6775_out0;
wire v_WENMULTI_5515_out0;
wire v_WENRAM_1134_out0;
wire v_WENRAM_2272_out0;
wire v_WEN_MULTI_1164_out0;
wire v_WEN_MULTI_5113_out0;
wire v_WRITE_EN_1582_out0;
wire v_W_EN_3377_out0;
wire v__0_out0;
wire v__1007_out0;
wire v__1008_out0;
wire v__1009_out0;
wire v__100_out0;
wire v__1010_out0;
wire v__1011_out0;
wire v__1012_out0;
wire v__1013_out0;
wire v__1014_out0;
wire v__1015_out0;
wire v__1016_out0;
wire v__1017_out0;
wire v__1018_out0;
wire v__1019_out0;
wire v__1020_out0;
wire v__1021_out0;
wire v__1022_out0;
wire v__1023_out0;
wire v__1048_out0;
wire v__1049_out0;
wire v__1050_out0;
wire v__1051_out0;
wire v__1052_out0;
wire v__1053_out0;
wire v__1054_out0;
wire v__1055_out0;
wire v__1056_out0;
wire v__1057_out0;
wire v__1058_out0;
wire v__1059_out0;
wire v__1060_out0;
wire v__1061_out0;
wire v__1062_out0;
wire v__1063_out0;
wire v__1064_out0;
wire v__1070_out0;
wire v__1071_out0;
wire v__1072_out0;
wire v__1073_out0;
wire v__1074_out0;
wire v__1075_out0;
wire v__1076_out0;
wire v__1077_out0;
wire v__1078_out0;
wire v__1079_out0;
wire v__1080_out0;
wire v__1081_out0;
wire v__1082_out0;
wire v__1083_out0;
wire v__1106_out0;
wire v__1109_out0;
wire v__1110_out0;
wire v__1111_out0;
wire v__1112_out0;
wire v__1113_out0;
wire v__1114_out0;
wire v__1115_out0;
wire v__1116_out0;
wire v__1117_out0;
wire v__1118_out0;
wire v__1119_out0;
wire v__1120_out0;
wire v__1121_out0;
wire v__1122_out0;
wire v__1123_out0;
wire v__1179_out0;
wire v__1180_out0;
wire v__1181_out0;
wire v__1185_out0;
wire v__1199_out0;
wire v__1203_out0;
wire v__1204_out0;
wire v__1220_out0;
wire v__1221_out0;
wire v__1222_out0;
wire v__1223_out0;
wire v__1224_out0;
wire v__1225_out0;
wire v__1226_out0;
wire v__1227_out0;
wire v__1228_out0;
wire v__1229_out0;
wire v__1230_out0;
wire v__1231_out0;
wire v__1232_out0;
wire v__1233_out0;
wire v__1234_out0;
wire v__1314_out0;
wire v__1331_out0;
wire v__1332_out0;
wire v__1333_out0;
wire v__1334_out0;
wire v__1335_out0;
wire v__1336_out0;
wire v__1337_out0;
wire v__1338_out0;
wire v__1339_out0;
wire v__1340_out0;
wire v__1341_out0;
wire v__1342_out0;
wire v__1343_out0;
wire v__1344_out0;
wire v__1345_out0;
wire v__1347_out0;
wire v__1348_out0;
wire v__1382_out0;
wire v__1382_out1;
wire v__1396_out0;
wire v__1401_out0;
wire v__1402_out0;
wire v__1403_out0;
wire v__1404_out0;
wire v__1407_out0;
wire v__142_out0;
wire v__1436_out0;
wire v__1443_out0;
wire v__1451_out0;
wire v__1456_out0;
wire v__1457_out0;
wire v__1458_out0;
wire v__1459_out0;
wire v__1460_out0;
wire v__1461_out0;
wire v__1462_out0;
wire v__1463_out0;
wire v__1464_out0;
wire v__1465_out0;
wire v__1466_out0;
wire v__1467_out0;
wire v__1468_out0;
wire v__1469_out0;
wire v__1470_out0;
wire v__1471_out0;
wire v__1488_out0;
wire v__1489_out0;
wire v__1490_out0;
wire v__1491_out0;
wire v__1492_out0;
wire v__1493_out0;
wire v__1494_out0;
wire v__1495_out0;
wire v__1496_out0;
wire v__1497_out0;
wire v__1498_out0;
wire v__1499_out0;
wire v__1500_out0;
wire v__1501_out0;
wire v__1502_out0;
wire v__1504_out0;
wire v__1505_out0;
wire v__1506_out0;
wire v__1507_out0;
wire v__1508_out0;
wire v__1509_out0;
wire v__1510_out0;
wire v__1511_out0;
wire v__1512_out0;
wire v__1513_out0;
wire v__1514_out0;
wire v__1515_out0;
wire v__1516_out0;
wire v__1517_out0;
wire v__1518_out0;
wire v__1521_out0;
wire v__1522_out0;
wire v__1523_out0;
wire v__1530_out0;
wire v__1531_out0;
wire v__1532_out0;
wire v__1533_out0;
wire v__1534_out0;
wire v__1535_out0;
wire v__1536_out0;
wire v__1537_out0;
wire v__1538_out0;
wire v__1539_out0;
wire v__1540_out0;
wire v__1541_out0;
wire v__1542_out0;
wire v__1543_out0;
wire v__1544_out0;
wire v__1550_out0;
wire v__1560_out0;
wire v__1576_out0;
wire v__1580_out0;
wire v__1581_out0;
wire v__1588_out0;
wire v__1590_out0;
wire v__1596_out0;
wire v__1597_out0;
wire v__159_out0;
wire v__160_out0;
wire v__163_out0;
wire v__164_out0;
wire v__1854_out0;
wire v__1863_out0;
wire v__1864_out0;
wire v__1865_out0;
wire v__1866_out0;
wire v__1867_out0;
wire v__1868_out0;
wire v__1869_out0;
wire v__1870_out0;
wire v__1871_out0;
wire v__1872_out0;
wire v__1873_out0;
wire v__1874_out0;
wire v__1875_out0;
wire v__1876_out0;
wire v__1877_out0;
wire v__1881_out0;
wire v__1882_out0;
wire v__1883_out0;
wire v__1884_out0;
wire v__1885_out0;
wire v__1886_out0;
wire v__1887_out0;
wire v__1888_out0;
wire v__1889_out0;
wire v__1890_out0;
wire v__1891_out0;
wire v__1892_out0;
wire v__1893_out0;
wire v__1894_out0;
wire v__1895_out0;
wire v__1905_out0;
wire v__1906_out0;
wire v__1907_out0;
wire v__1908_out0;
wire v__1909_out0;
wire v__1910_out0;
wire v__1911_out0;
wire v__1912_out0;
wire v__1913_out0;
wire v__1914_out0;
wire v__1915_out0;
wire v__1916_out0;
wire v__1917_out0;
wire v__1918_out0;
wire v__1919_out0;
wire v__1920_out0;
wire v__1933_out0;
wire v__1934_out0;
wire v__1935_out0;
wire v__1936_out0;
wire v__1937_out0;
wire v__1938_out0;
wire v__1939_out0;
wire v__1940_out0;
wire v__1941_out0;
wire v__1942_out0;
wire v__1943_out0;
wire v__1944_out0;
wire v__1945_out0;
wire v__1946_out0;
wire v__1947_out0;
wire v__1_out0;
wire v__201_out0;
wire v__212_out0;
wire v__21_out0;
wire v__2211_out1;
wire v__2244_out0;
wire v__2245_out0;
wire v__2248_out0;
wire v__2248_out1;
wire v__2251_out0;
wire v__229_out0;
wire v__2300_out0;
wire v__2301_out0;
wire v__230_out0;
wire v__231_out0;
wire v__232_out0;
wire v__233_out0;
wire v__234_out0;
wire v__2350_out0;
wire v__2351_out0;
wire v__2358_out1;
wire v__2359_out0;
wire v__235_out0;
wire v__2361_out0;
wire v__236_out0;
wire v__2370_out0;
wire v__237_out0;
wire v__238_out0;
wire v__239_out0;
wire v__240_out0;
wire v__241_out0;
wire v__242_out0;
wire v__243_out0;
wire v__246_out0;
wire v__247_out0;
wire v__248_out0;
wire v__249_out0;
wire v__250_out0;
wire v__251_out0;
wire v__252_out0;
wire v__253_out0;
wire v__254_out0;
wire v__255_out0;
wire v__256_out0;
wire v__257_out0;
wire v__258_out0;
wire v__259_out0;
wire v__260_out0;
wire v__277_out0;
wire v__278_out0;
wire v__279_out0;
wire v__280_out0;
wire v__281_out0;
wire v__282_out0;
wire v__283_out0;
wire v__284_out0;
wire v__2859_out0;
wire v__2859_out1;
wire v__285_out0;
wire v__286_out0;
wire v__2870_out0;
wire v__2870_out1;
wire v__287_out0;
wire v__288_out0;
wire v__289_out0;
wire v__290_out0;
wire v__291_out0;
wire v__31_out0;
wire v__3340_out0;
wire v__3341_out0;
wire v__3342_out0;
wire v__3343_out0;
wire v__3344_out0;
wire v__3345_out0;
wire v__3346_out0;
wire v__3347_out0;
wire v__3348_out0;
wire v__3349_out0;
wire v__3350_out0;
wire v__3351_out0;
wire v__3352_out0;
wire v__3353_out0;
wire v__3354_out0;
wire v__3355_out0;
wire v__3356_out0;
wire v__3357_out0;
wire v__3358_out0;
wire v__3359_out0;
wire v__3360_out0;
wire v__3361_out0;
wire v__3362_out0;
wire v__3363_out0;
wire v__3364_out0;
wire v__3365_out0;
wire v__3366_out0;
wire v__3367_out0;
wire v__3368_out0;
wire v__3369_out0;
wire v__3376_out0;
wire v__3376_out1;
wire v__3467_out1;
wire v__3471_out0;
wire v__3482_out0;
wire v__3487_out0;
wire v__3756_out0;
wire v__3757_out0;
wire v__3758_out0;
wire v__3759_out0;
wire v__3760_out0;
wire v__3761_out0;
wire v__3762_out0;
wire v__3763_out0;
wire v__3764_out0;
wire v__3765_out0;
wire v__3766_out0;
wire v__3767_out0;
wire v__3768_out0;
wire v__3769_out0;
wire v__3770_out0;
wire v__40_out0;
wire v__41_out0;
wire v__4282_out0;
wire v__4283_out0;
wire v__4284_out0;
wire v__4285_out0;
wire v__4286_out0;
wire v__4287_out0;
wire v__4288_out0;
wire v__4289_out0;
wire v__4290_out0;
wire v__4291_out0;
wire v__4292_out0;
wire v__4293_out0;
wire v__4294_out0;
wire v__4295_out0;
wire v__4296_out0;
wire v__4305_out0;
wire v__4306_out0;
wire v__4315_out0;
wire v__4316_out0;
wire v__4317_out0;
wire v__4318_out0;
wire v__4319_out0;
wire v__4320_out0;
wire v__4321_out0;
wire v__4322_out0;
wire v__4323_out0;
wire v__4324_out0;
wire v__4325_out0;
wire v__4326_out0;
wire v__4327_out0;
wire v__4328_out0;
wire v__4329_out0;
wire v__4343_out0;
wire v__4344_out0;
wire v__4345_out0;
wire v__4353_out0;
wire v__4354_out0;
wire v__5111_out0;
wire v__5112_out0;
wire v__5115_out0;
wire v__5116_out0;
wire v__5127_out0;
wire v__5128_out0;
wire v__5129_out0;
wire v__5130_out0;
wire v__5131_out0;
wire v__5132_out0;
wire v__5133_out0;
wire v__5134_out0;
wire v__5135_out0;
wire v__5136_out0;
wire v__5137_out0;
wire v__5138_out0;
wire v__5139_out0;
wire v__5140_out0;
wire v__5141_out0;
wire v__5157_out0;
wire v__5160_out0;
wire v__5164_out1;
wire v__5184_out0;
wire v__5185_out0;
wire v__5264_out0;
wire v__5265_out0;
wire v__5275_out0;
wire v__5276_out0;
wire v__5277_out0;
wire v__5278_out0;
wire v__5279_out0;
wire v__5280_out0;
wire v__5281_out0;
wire v__5282_out0;
wire v__5283_out0;
wire v__5284_out0;
wire v__5285_out0;
wire v__5286_out0;
wire v__5287_out0;
wire v__5288_out0;
wire v__5289_out0;
wire v__5290_out0;
wire v__5304_out0;
wire v__5305_out0;
wire v__5308_out0;
wire v__5317_out0;
wire v__5324_out0;
wire v__5343_out0;
wire v__5344_out0;
wire v__5347_out1;
wire v__5349_out0;
wire v__5350_out0;
wire v__5351_out0;
wire v__5352_out0;
wire v__5353_out0;
wire v__5354_out0;
wire v__5355_out0;
wire v__5356_out0;
wire v__5357_out0;
wire v__5358_out0;
wire v__5359_out0;
wire v__5360_out0;
wire v__5361_out0;
wire v__5362_out0;
wire v__5363_out0;
wire v__5367_out0;
wire v__5414_out0;
wire v__5415_out0;
wire v__5416_out0;
wire v__5417_out0;
wire v__5418_out0;
wire v__5419_out0;
wire v__5420_out0;
wire v__5421_out0;
wire v__5422_out0;
wire v__5423_out0;
wire v__5424_out0;
wire v__5425_out0;
wire v__5426_out0;
wire v__5427_out0;
wire v__5428_out0;
wire v__5463_out0;
wire v__5464_out0;
wire v__5465_out0;
wire v__5466_out0;
wire v__5467_out0;
wire v__5468_out0;
wire v__5469_out0;
wire v__5470_out0;
wire v__5471_out0;
wire v__5472_out0;
wire v__5473_out0;
wire v__5474_out0;
wire v__5475_out0;
wire v__5476_out0;
wire v__5477_out0;
wire v__5487_out0;
wire v__5488_out0;
wire v__5518_out0;
wire v__5532_out0;
wire v__5559_out1;
wire v__577_out0;
wire v__584_out0;
wire v__6535_out0;
wire v__6593_out0;
wire v__6594_out0;
wire v__6597_out0;
wire v__6599_out0;
wire v__6600_out0;
wire v__6601_out0;
wire v__6602_out0;
wire v__6603_out0;
wire v__6604_out0;
wire v__6605_out0;
wire v__6606_out0;
wire v__6607_out0;
wire v__6608_out0;
wire v__6609_out0;
wire v__6610_out0;
wire v__6611_out0;
wire v__6612_out0;
wire v__6613_out0;
wire v__6614_out0;
wire v__6618_out0;
wire v__6624_out0;
wire v__6625_out0;
wire v__6626_out0;
wire v__6627_out0;
wire v__6628_out0;
wire v__6629_out0;
wire v__6630_out0;
wire v__6631_out0;
wire v__6632_out0;
wire v__6633_out0;
wire v__6634_out0;
wire v__6635_out0;
wire v__6636_out0;
wire v__6637_out0;
wire v__6638_out0;
wire v__6659_out0;
wire v__6660_out0;
wire v__6679_out0;
wire v__6680_out0;
wire v__6683_out0;
wire v__6703_out0;
wire v__6714_out0;
wire v__6715_out0;
wire v__6756_out0;
wire v__6757_out0;
wire v__6758_out0;
wire v__6759_out0;
wire v__6760_out0;
wire v__6761_out0;
wire v__6762_out0;
wire v__6763_out0;
wire v__6764_out0;
wire v__6765_out0;
wire v__6766_out0;
wire v__6767_out0;
wire v__6768_out0;
wire v__6769_out0;
wire v__6770_out0;
wire v__831_out0;
wire v__832_out0;
wire v__844_out0;
wire v__845_out0;
wire v__846_out0;
wire v__853_out0;
wire v__854_out0;
wire v__867_out0;
wire v__868_out0;
wire v__869_out0;
wire v__870_out0;
wire v__871_out0;
wire v__872_out0;
wire v__873_out0;
wire v__874_out0;
wire v__875_out0;
wire v__876_out0;
wire v__877_out0;
wire v__878_out0;
wire v__879_out0;
wire v__880_out0;
wire v__881_out0;
wire v__88_out0;
wire v__917_out0;
wire v__926_out0;
wire v__927_out0;
wire v__92_out0;
wire v__931_out0;
wire v__94_out0;
wire v__965_out0;
wire v__966_out0;
wire v__967_out0;
wire v__968_out0;
wire v__969_out0;
wire v__970_out0;
wire v__971_out0;
wire v__972_out0;
wire v__973_out0;
wire v__974_out0;
wire v__975_out0;
wire v__976_out0;
wire v__977_out0;
wire v__978_out0;
wire v__979_out0;
wire v__97_out0;
wire v__986_out0;
wire v__98_out0;
wire v_done_receiving_5219_out0;
wire v_transmit_INSTRUCTION_1304_out0;
wire v_tx_Overflow_1349_out0;
wire v_tx_in_progress_1449_out0;
wire v_tx_in_progress_1925_out0;
wire v_uart_5478_out0;

always @(posedge clk) v_FF1_26_out0 <= v_BYTE_READY_1393_out0;
always @(posedge clk) v_FF2_43_out0 <= v__2248_out1;
always @(posedge clk) v_FF6_58_out0 <= v_ENABLE_1292_out0 ? v_MUX5_6574_out0 : v_FF6_58_out0;
always @(posedge clk) v_REG1_210_out0 <= v_G12_5202_out0 ? v_MUX4_1295_out0 : v_REG1_210_out0;
v_ROM1_225 I1 (v_ROM1_225_out0, v_REG1_3500_out0, clk);
always @(posedge clk) v_FF4_226_out0 <= v_ENABLE_1292_out0 ? v_MUX3_3503_out0 : v_FF4_226_out0;
v_RAM1_930 I1 (v_RAM1_930_out0, v_MUX3_1571_out0, v_MUX2_1561_out0, v_G1_5271_out0, clk);
always @(posedge clk) v_FF1_956_out0 <= v_ENABLE_1292_out0 ? v_SEL1_6622_out0 : v_FF1_956_out0;
always @(posedge clk) v_IHOLD_REGISTER_983_out0 <= v_NORMAL_93_out0 ? v_RAM_OUT_855_out0 : v_IHOLD_REGISTER_983_out0;
always @(posedge clk) v_REG1_1128_out0 <= v_D1_4350_out1 ? v_DIN3_5083_out0 : v_REG1_1128_out0;
always @(posedge clk) v_FF7_1302_out0 <= v_G24_5196_out0;
always @(posedge clk) v_FF7_1303_out0 <= v_G24_5197_out0;
always @(posedge clk) v_REG1_1306_out0 <= v_ENABLE_859_out0 ? v__1482_out0 : v_REG1_1306_out0;
always @(posedge clk) v_FF2_1362_out0 <= v_INSTRUCTION_32_out0 ? v_G3_5370_out0 : v_FF2_1362_out0;
always @(posedge clk) v_FF2_1383_out0 <= v_ENABLE_1292_out0 ? v_MUX1_1279_out0 : v_FF2_1383_out0;
always @(posedge clk) v_FF1_2303_out0 <= v_EN_1423_out0 ? v_G1_1318_out0 : v_FF1_2303_out0;
always @(posedge clk) v_FF1_2304_out0 <= v_EN_1424_out0 ? v_G1_1319_out0 : v_FF1_2304_out0;
always @(posedge clk) v_FF1_2305_out0 <= v_EN_1425_out0 ? v_G1_1320_out0 : v_FF1_2305_out0;
always @(posedge clk) v_FF1_2306_out0 <= v_EN_1426_out0 ? v_G1_1321_out0 : v_FF1_2306_out0;
always @(posedge clk) v_FF1_2307_out0 <= v_EN_1427_out0 ? v_G1_1322_out0 : v_FF1_2307_out0;
always @(posedge clk) v_FF1_2308_out0 <= v_EN_1428_out0 ? v_G1_1323_out0 : v_FF1_2308_out0;
always @(posedge clk) v_FF1_2309_out0 <= v_EN_1429_out0 ? v_G1_1324_out0 : v_FF1_2309_out0;
always @(posedge clk) v_FF1_2310_out0 <= v_EN_1430_out0 ? v_G1_1325_out0 : v_FF1_2310_out0;
always @(posedge clk) v_REG3_2317_out0 <= v_D1_4350_out3 ? v_DIN3_5083_out0 : v_REG3_2317_out0;
always @(posedge clk) v_FF7_2334_out0 <= v_ENABLE_1292_out0 ? v_MUX6_5401_out0 : v_FF7_2334_out0;
always @(posedge clk) v_FF5_3484_out0 <= v_ENABLE_1292_out0 ? v_MUX4_1568_out0 : v_FF5_3484_out0;
always @(posedge clk) v_REG1_3500_out0 <= v_EQ3_2871_out0 ? v_A1_5433_out0 : v_REG1_3500_out0;
always @(posedge clk) v_FF9_4333_out0 <= v_ENABLE_1292_out0 ? v_MUX8_1316_out0 : v_FF9_4333_out0;
always @(posedge clk) v_FF1_5090_out0 <= v_G3_1435_out0 ? v_G2_5313_out0 : v_FF1_5090_out0;
always @(posedge clk) v_REG1_5108_out0 <= v__261_out0;
always @(posedge clk) v_FF3_5175_out0 <= v_G8_6721_out0;
always @(posedge clk) v_REG1_5190_out0 <= v_G8_9_out0 ? v_OUT_1480_out0 : v_REG1_5190_out0;
always @(posedge clk) v_FF8_5337_out0 <= v_G21_1856_out0;
always @(posedge clk) v_FF8_5338_out0 <= v_G21_1857_out0;
always @(posedge clk) v_REG0_5368_out0 <= v_D1_4350_out0 ? v_DIN3_5083_out0 : v_REG0_5368_out0;
always @(posedge clk) v_FF3_5435_out0 <= v_ENABLE_1292_out0 ? v_MUX2_2175_out0 : v_FF3_5435_out0;
always @(posedge clk) v_FF1_5442_out0 <= v__2248_out0;
always @(posedge clk) v_FF2_5444_out0 <= v_FF1_6658_out0;
always @(posedge clk) v_REG1_5479_out0 <= v_G2_3380_out0 ? v_COUT_1898_out0 : v_REG1_5479_out0;
always @(posedge clk) v_FF8_5523_out0 <= v_ENABLE_1292_out0 ? v_MUX7_5145_out0 : v_FF8_5523_out0;
always @(posedge clk) v_REG2_6035_out0 <= v_D1_4350_out2 ? v_DIN3_5083_out0 : v_REG2_6035_out0;
always @(posedge clk) v_REG1_6571_out0 <= v_COUT_5377_out0;
always @(posedge clk) v_FF1_6658_out0 <= v_ROM1_225_out0;
assign v_C11_6781_out0 = 6'h0;
assign v_C1_6623_out0 = 8'h0;
assign v_C1_6547_out0 = 8'h0;
assign v_C5_6541_out0 = 1'h1;
assign v_C1_5558_out0 = 2'h0;
assign v_C10_5536_out0 = 5'h1f;
assign v_C9_5492_out0 = 6'h3f;
assign v_C14_5312_out0 = 5'h1;
assign v_C1_5309_out0 = 1'h0;
assign v_C2_5297_out0 = 12'h7ff;
assign v_C4_5227_out0 = 1'h1;
assign v_C6_5086_out0 = 1'h1;
assign v_C1_5085_out0 = 5'h0;
assign v_C1_5084_out0 = 5'h0;
assign v_C1_5082_out0 = 4'h0;
assign v_C1_5063_out0 = 8'h0;
assign v_C1_5058_out0 = 1'h0;
assign v_C1_4338_out0 = 1'h0;
assign v_2_3472_out0 = 1'h1;
assign v_C1_3397_out0 = 4'h0;
assign v_C1_3337_out0 = 2'h0;
assign v_C3_2314_out0 = 1'h0;
assign v_C11_2218_out0 = 16'hffff;
assign v_C1_1564_out0 = 12'h0;
assign v_C1_1562_out0 = 2'h0;
assign v_C9_1477_out0 = 1'h0;
assign v_C8_1346_out0 = 5'h0;
assign v_C5_1312_out0 = 16'hffff;
assign v_C4_1264_out0 = 5'h0;
assign v_C1_1182_out0 = 12'h7f6;
assign v_C2_1176_out0 = 12'h0;
assign v_C7_1108_out0 = 1'h0;
assign v_C13_1065_out0 = 16'h0;
assign v_C12_1029_out0 = 6'hf;
assign v_C1_980_out0 = 4'h4;
assign v_C7_912_out0 = 16'h0;
assign v_C10_888_out0 = 1'h1;
assign v_C_883_out0 = 12'h1;
assign v_C15_847_out0 = 16'hffff;
assign v_C14_822_out0 = 1'h1;
assign v_C12_565_out0 = 1'h1;
assign v_C1_294_out0 = 11'h0;
assign v_C1_293_out0 = 1'h0;
assign v_C1_211_out0 = 1'h1;
assign v_C13_196_out0 = 6'h31;
assign v_ROR_34_out0 = 2'h3;
assign v_Q_144_out0 = v_FF1_2303_out0;
assign v_Q_145_out0 = v_FF1_2304_out0;
assign v_Q_146_out0 = v_FF1_2305_out0;
assign v_Q_147_out0 = v_FF1_2306_out0;
assign v_Q_148_out0 = v_FF1_2307_out0;
assign v_Q_149_out0 = v_FF1_2308_out0;
assign v_Q_150_out0 = v_FF1_2309_out0;
assign v_Q_151_out0 = v_FF1_2310_out0;
assign v_EQ4_560_out0 = v_REG1_3500_out0 == 12'h0;
assign v_R0_828_out0 = v_REG0_5368_out0;
assign v_Q6_924_out0 = v_FF7_1302_out0;
assign v_Q6_925_out0 = v_FF7_1303_out0;
assign v_IR_1380_out0 = v_IHOLD_REGISTER_983_out0;
assign v__1406_out0 = { v_FF1_5442_out0,v_FF2_43_out0 };
assign v__1443_out0 = v_REG1_1306_out0[0:0];
assign v__1443_out1 = v_REG1_1306_out0[7:7];
assign v_OUT_1480_out0 = v_REG1_1306_out0;
assign v_R2_1484_out0 = v_REG2_6035_out0;
assign v_C_1559_out0 = v_REG1_5479_out0;
assign v_C_1563_out0 = v_REG1_5479_out0;
assign v_EN_2191_out0 = v_C5_6541_out0;
assign v_R3_2273_out0 = v_REG3_2317_out0;
assign v__2870_out0 = v_REG1_5108_out0[0:0];
assign v__2870_out1 = v_REG1_5108_out0[1:1];
assign v_Q7_3382_out0 = v_FF8_5337_out0;
assign v_Q7_3383_out0 = v_FF8_5338_out0;
assign v_NEG1_3398_out0 = v_C9_5492_out0;
assign v__3490_out0 = v_IHOLD_REGISTER_983_out0[11:0];
assign v__3490_out1 = v_IHOLD_REGISTER_983_out0[15:4];
assign v_RAM_OUT_3506_out0 = v_RAM1_930_out0;
assign v_RECEIVERSTREAM_3751_out0 = v_REG1_5190_out0;
assign v_Q_3786_out0 = v_FF3_5175_out0;
assign v_TRANSMITER_OVERFLOW_4268_out0 = v_FF2_1362_out0;
assign v_R1_4311_out0 = v_REG1_1128_out0;
assign v_0B00001_5193_out0 = v_C14_5312_out0;
assign v_Q_5226_out0 = v_REG1_5108_out0;
assign v_0_5269_out0 = v_C7_1108_out0;
assign v_G2_5313_out0 = ! v_FF1_5090_out0;
assign v_A_5323_out0 = v_C_883_out0;
assign {v_A1_5433_out1,v_A1_5433_out0 } = v_C2_1176_out0 + v_REG1_3500_out0 + v_C1_211_out0;
assign v_DIV_INSTRUCTION_5560_out0 = v_DIV_INST_1133_out0;
assign v_FLOAT_INST16_6621_out0 = v_FF1_5090_out0;
assign v__31_out0 = v_A_5323_out0[10:10];
assign v__88_out0 = v_A_5323_out0[7:7];
assign v__92_out0 = v_A_5323_out0[3:3];
assign v__142_out0 = v_A_5323_out0[2:2];
assign v_RECEIVER_STREAM_276_out0 = v_RECEIVERSTREAM_3751_out0;
assign v_Q_566_out0 = v__1406_out0;
assign v_G5_587_out0 = ! v_EN_2191_out0;
assign v_Q2_823_out0 = v_Q_144_out0;
assign v_Q2_824_out0 = v_Q_148_out0;
assign v_RAM_OUT_855_out0 = v_RAM_OUT_3506_out0;
assign v__917_out0 = v_A_5323_out0[11:11];
assign v_G10_950_out0 = !(v_Q_145_out0 || v_Q_144_out0);
assign v_G10_951_out0 = !(v_Q_149_out0 || v_Q_148_out0);
assign v_G4_958_out0 = v_Q_147_out0 && v_Q_145_out0;
assign v_G4_959_out0 = v_Q_151_out0 && v_Q_149_out0;
assign v__986_out0 = v_A_5323_out0[5:5];
assign v_G28_1025_out0 = v_Q7_3382_out0 && v_Q6_924_out0;
assign v_G28_1026_out0 = v_Q7_3383_out0 && v_Q6_925_out0;
assign v_Q1_1028_out0 = v__2870_out1;
assign v__1106_out0 = v_A_5323_out0[8:8];
assign v_EQ10_1131_out0 = v__3490_out1 == 4'h3;
assign v_TX_OVERFLOW_1184_out0 = v_TRANSMITER_OVERFLOW_4268_out0;
assign v_COUT_1330_out0 = v_A1_5433_out1;
assign v_R3TEST_1400_out0 = v_R3_2273_out0;
assign v_G2_1452_out0 = ((v_Q_147_out0 && !v_Q_145_out0) || (!v_Q_147_out0) && v_Q_145_out0);
assign v_G2_1453_out0 = ((v_Q_151_out0 && !v_Q_149_out0) || (!v_Q_151_out0) && v_Q_149_out0);
assign v__1523_out0 = v_A_5323_out0[1:1];
assign v_R0TEST_1552_out0 = v_R0_828_out0;
assign v__1590_out0 = v_A_5323_out0[4:4];
assign v_NOTUSED_2250_out0 = v__1443_out0;
assign v_G23_2368_out0 = ! v_Q7_3382_out0;
assign v_G23_2369_out0 = ! v_Q7_3383_out0;
assign v_EQ3_2871_out0 = v_Q_5226_out0 == 2'h3;
assign v_IR_3489_out0 = v_IR_1380_out0;
assign v__3525_out0 = { v_Q7_3382_out0,v_Q6_924_out0 };
assign v__3526_out0 = { v_Q7_3383_out0,v_Q6_925_out0 };
assign v_C_4256_out0 = v_C_1563_out0;
assign v_G1_4279_out0 = ! v_Q_147_out0;
assign v_G1_4280_out0 = ! v_Q_151_out0;
assign v_Q3_4301_out0 = v_Q_146_out0;
assign v_Q3_4302_out0 = v_Q_150_out0;
assign v_Q1_4358_out0 = v_Q_145_out0;
assign v_Q1_4359_out0 = v_Q_149_out0;
assign v_G9_5075_out0 = v_Q_147_out0 && v_Q_146_out0;
assign v_G9_5076_out0 = v_Q_151_out0 && v_Q_150_out0;
assign v_FLOATING_INSTRUCTION_5118_out0 = v_FLOAT_INST16_6621_out0;
assign v_R1TEST_5162_out0 = v_R1_4311_out0;
assign v_G24_5196_out0 = ((v_Q7_3382_out0 && !v_Q6_924_out0) || (!v_Q7_3382_out0) && v_Q6_924_out0);
assign v_G24_5197_out0 = ((v_Q7_3383_out0 && !v_Q6_925_out0) || (!v_Q7_3383_out0) && v_Q6_925_out0);
assign v_R2TEST_5270_out0 = v_R2_1484_out0;
assign v_Q0_5512_out0 = v_Q_147_out0;
assign v_Q0_5513_out0 = v_Q_151_out0;
assign v_RAM_OUT_5521_out0 = v_RAM_OUT_3506_out0;
assign v__5532_out0 = v_A_5323_out0[9:9];
assign v_Q0_6576_out0 = v__2870_out0;
assign v__6599_out0 = v_A_5323_out0[6:6];
assign v_NOUSED_6647_out0 = v__3490_out0;
assign v__6683_out0 = v_A_5323_out0[0:0];
assign v_DIV_INSTRUCTION_6717_out0 = v_DIV_INSTRUCTION_5560_out0;
assign v_EQ2_5_out0 = v_Q_566_out0 == 2'h2;
assign v_R3TEST_61_out0 = v_R3TEST_1400_out0;
assign v__112_out0 = v_RAM_OUT_855_out0[11:0];
assign v__112_out1 = v_RAM_OUT_855_out0[15:4];
assign v_4BITCOUNTER_157_out0 = v__3525_out0;
assign v_4BITCOUNTER_158_out0 = v__3526_out0;
assign v_RAM_OUT_200_out0 = v_RAM_OUT_5521_out0;
assign v_EQ4_296_out0 = v_Q_566_out0 == 2'h0;
assign v_G6_569_out0 = v_G4_958_out0 && v_Q_144_out0;
assign v_G6_570_out0 = v_G4_959_out0 && v_Q_148_out0;
assign v_IR_915_out0 = v_IR_3489_out0;
assign v_G12_1107_out0 = ! v_Q1_1028_out0;
assign v_EQ1_1238_out0 = v_Q_566_out0 == 2'h1;
assign v_DIV_INSTRUCTION_1602_out0 = v_DIV_INSTRUCTION_6717_out0;
assign v_G3_1625_out0 = v_G5_587_out0 && v_Q1_1028_out0;
assign v_G38_1903_out0 = v_Q2_823_out0 || v_Q3_4301_out0;
assign v_G38_1904_out0 = v_Q2_824_out0 || v_Q3_4302_out0;
assign v_Q0_2184_out0 = v_Q0_5512_out0;
assign v_Q0_2185_out0 = v_Q0_5513_out0;
assign v_C_2366_out0 = v_C_4256_out0;
assign v__2859_out0 = v_Q_566_out0[0:0];
assign v__2859_out1 = v_Q_566_out0[1:1];
assign v_Q2_3378_out0 = v_Q2_823_out0;
assign v_Q2_3379_out0 = v_Q2_824_out0;
assign v_G3_3385_out0 = ((v_G4_958_out0 && !v_Q_144_out0) || (!v_G4_958_out0) && v_Q_144_out0);
assign v_G3_3386_out0 = ((v_G4_959_out0 && !v_Q_148_out0) || (!v_G4_959_out0) && v_Q_148_out0);
assign v_G37_3388_out0 = v_Q1_4358_out0 || v_Q0_5512_out0;
assign v_G37_3389_out0 = v_Q1_4359_out0 || v_Q0_5513_out0;
assign v_Q1_3390_out0 = v_Q1_4358_out0;
assign v_Q1_3391_out0 = v_Q1_4359_out0;
assign v_G4_3394_out0 = ! v_Q0_6576_out0;
assign v_R0TEST_3439_out0 = v_R0TEST_1552_out0;
assign v_D_3774_out0 = v_G2_1452_out0;
assign v_D_3776_out0 = v_G1_4279_out0;
assign v_D_3778_out0 = v_G2_1453_out0;
assign v_D_3780_out0 = v_G1_4280_out0;
assign v_G11_4258_out0 = v_EN_2191_out0 && v_Q0_6576_out0;
assign v_G2_5068_out0 = ! v_EQ3_2871_out0;
assign v_EN_5147_out0 = v_G28_1025_out0;
assign v_EN_5148_out0 = v_G28_1026_out0;
assign v_R1TEST_5168_out0 = v_R1TEST_5162_out0;
assign v_Q3_5177_out0 = v_Q3_4301_out0;
assign v_Q3_5178_out0 = v_Q3_4302_out0;
assign v_RECEIVER_stream_5189_out0 = v_RECEIVER_STREAM_276_out0;
assign v_G8_5222_out0 = !(v_G9_5075_out0 && v_G10_950_out0);
assign v_G8_5223_out0 = !(v_G9_5076_out0 && v_G10_951_out0);
assign v_G1_5318_out0 = ((v_EN_2191_out0 && !v_Q0_6576_out0) || (!v_EN_2191_out0) && v_Q0_6576_out0);
assign v_G22_5405_out0 = v_G23_2368_out0 && v_Q6_924_out0;
assign v_G22_5406_out0 = v_G23_2369_out0 && v_Q6_925_out0;
assign v_R2TEST_5407_out0 = v_R2TEST_5270_out0;
assign v_SHIFHT_ENABLE_6652_out0 = v_G28_1025_out0;
assign v_SHIFHT_ENABLE_6653_out0 = v_G28_1026_out0;
assign v_EQ3_6655_out0 = v_Q_566_out0 == 2'h3;
assign v_FLOATING_INS_6796_out0 = v_FLOATING_INSTRUCTION_5118_out0;
assign v_4BITCOUNTER_4_out0 = v_4BITCOUNTER_158_out0;
assign v_EQ6_11_out0 = v_4BITCOUNTER_157_out0 == 2'h2;
assign v_R3_38_out0 = v_R3TEST_61_out0;
assign v_NORMAL_93_out0 = v_EQ1_1238_out0;
assign v_Q1_152_out0 = v__2859_out1;
assign v_EQ1_156_out0 = v__112_out1 == 4'h0;
assign v_EXEC1LS_209_out0 = v_EQ2_5_out0;
assign v_Q0_303_out0 = v__2859_out0;
assign v_G7_586_out0 = v_G11_4258_out0 && v_G12_1107_out0;
assign v_9_834_out0 = v_G8_5222_out0;
assign v_9_835_out0 = v_G8_5223_out0;
assign v_FLAOTING_INSTRUCTION_908_out0 = v_FLOATING_INS_6796_out0;
assign v_EQ6_961_out0 = v__112_out1 == 4'h5;
assign v_R1_1003_out0 = v_R1TEST_5168_out0;
assign v_EQ9_1165_out0 = v__112_out1 == 4'h3;
assign v_EQ8_1194_out0 = v__112_out1 == 4'h7;
assign v_EQ11_1196_out0 = v__112_out1 == 4'h1;
assign v_ADRESS_1239_out0 = v__112_out0;
assign v_G5_1260_out0 = ((v_G6_569_out0 && !v_Q_146_out0) || (!v_G6_569_out0) && v_Q_146_out0);
assign v_G5_1261_out0 = ((v_G6_570_out0 && !v_Q_150_out0) || (!v_G6_570_out0) && v_Q_150_out0);
assign v_R0_1392_out0 = v_R0TEST_3439_out0;
assign v_IR_1413_out0 = v_IR_915_out0;
assign v_G1_1418_out0 = v_EQ4_560_out0 && v_G2_5068_out0;
assign v_EN_1423_out0 = v_EN_5147_out0;
assign v_EN_1424_out0 = v_EN_5147_out0;
assign v_EN_1425_out0 = v_EN_5147_out0;
assign v_EN_1426_out0 = v_EN_5147_out0;
assign v_EN_1427_out0 = v_EN_5148_out0;
assign v_EN_1428_out0 = v_EN_5148_out0;
assign v_EN_1429_out0 = v_EN_5148_out0;
assign v_EN_1430_out0 = v_EN_5148_out0;
assign v_START_1476_out0 = v_EQ4_296_out0;
assign v_G36_1528_out0 = !(v_G38_1903_out0 || v_G37_3388_out0);
assign v_G36_1529_out0 = !(v_G38_1904_out0 || v_G37_3389_out0);
assign v_EXEC2LS_1554_out0 = v_EQ3_6655_out0;
assign v_EQ7_1608_out0 = v__112_out1 == 4'h6;
assign v_DIV_INSTRUCTION_2254_out0 = v_DIV_INSTRUCTION_1602_out0;
assign v_4BITCOUNTER_2360_out0 = v_4BITCOUNTER_157_out0;
assign v_EQ5_2372_out0 = v__112_out1 == 4'h4;
assign v__3476_out0 = { v_RECEIVER_stream_5189_out0,v_C1_6547_out0 };
assign v_EQ3_3505_out0 = v__112_out1 == 4'h2;
assign v_D_3773_out0 = v_G3_3385_out0;
assign v_D_3777_out0 = v_G3_3386_out0;
assign v_SHIFT_ENABLE_4275_out0 = v_SHIFHT_ENABLE_6652_out0;
assign v_EQ5_4313_out0 = v_4BITCOUNTER_157_out0 == 2'h0;
assign v__4824_out0 = { v_C1_6547_out0,v_RECEIVER_stream_5189_out0 };
assign v_EQ2_4827_out0 = v_4BITCOUNTER_157_out0 == 2'h1;
assign v__5073_out0 = { v_Q0_2184_out0,v_Q1_3390_out0 };
assign v__5074_out0 = { v_Q0_2185_out0,v_Q1_3391_out0 };
assign v_G10_5272_out0 = v_G4_3394_out0 && v_Q1_1028_out0;
assign v_R2_5364_out0 = v_R2TEST_5407_out0;
assign v_EQ2_5404_out0 = v_4BITCOUNTER_158_out0 == 2'h0;
assign v_RESET_5499_out0 = v_G8_5222_out0;
assign v_RESET_5500_out0 = v_G8_5222_out0;
assign v_RESET_5501_out0 = v_G8_5222_out0;
assign v_RESET_5502_out0 = v_G8_5222_out0;
assign v_RESET_5503_out0 = v_G8_5223_out0;
assign v_RESET_5504_out0 = v_G8_5223_out0;
assign v_RESET_5505_out0 = v_G8_5223_out0;
assign v_RESET_5506_out0 = v_G8_5223_out0;
assign v_RAM_OUT_5519_out0 = v_RAM_OUT_200_out0;
assign v_RECEIVER_STREAM_6544_out0 = v_RECEIVER_stream_5189_out0;
assign v__2_out0 = v_IR_1413_out0[14:12];
assign v_R3_20_out0 = v_R3_38_out0;
assign v_MUX1_314_out0 = v_G1_1418_out0 ? v_C4_5227_out0 : v_FF2_5444_out0;
assign v_G1_573_out0 = ! v_Q0_303_out0;
assign v_G3_843_out0 = ! v_FLAOTING_INSTRUCTION_908_out0;
assign v_JMI_948_out0 = v_EQ6_961_out0;
assign v_ADRESS_1141_out0 = v_ADRESS_1239_out0;
assign v_R0_1237_out0 = v_R0_1392_out0;
assign v__1267_out0 = v_IR_1413_out0[1:0];
assign v_R1_1282_out0 = v_R1_1003_out0;
assign v_G2_1293_out0 = v_EQ9_1165_out0 || v_EQ10_1131_out0;
assign v_G1_1318_out0 = v_RESET_5499_out0 && v_D_3773_out0;
assign v_G1_1319_out0 = v_RESET_5500_out0 && v_D_3774_out0;
assign v_G1_1321_out0 = v_RESET_5502_out0 && v_D_3776_out0;
assign v_G1_1322_out0 = v_RESET_5503_out0 && v_D_3777_out0;
assign v_G1_1323_out0 = v_RESET_5504_out0 && v_D_3778_out0;
assign v_G1_1325_out0 = v_RESET_5506_out0 && v_D_3780_out0;
assign v_4BITCOUNTER_1419_out0 = v_4BITCOUNTER_2360_out0;
assign v__1444_out0 = { v__5073_out0,v_Q2_3378_out0 };
assign v__1445_out0 = { v__5074_out0,v_Q2_3379_out0 };
assign v_G6_2214_out0 = v_G10_5272_out0 || v_G3_1625_out0;
assign v_FLOAT_2247_out0 = v_EQ3_3505_out0;
assign v_RECEIVE_REGISTER_2841_out0 = v_RECEIVER_STREAM_6544_out0;
assign v_G2_3336_out0 = ! v_Q1_152_out0;
assign v_EXEC1LS_3338_out0 = v_EXEC1LS_209_out0;
assign v_G13_3477_out0 = v_Q0_303_out0 && v_Q1_152_out0;
assign v__3482_out0 = v_IR_1413_out0[15:15];
assign v_D_3775_out0 = v_G5_1260_out0;
assign v_D_3779_out0 = v_G5_1261_out0;
assign v_JMP_4342_out0 = v_EQ5_2372_out0;
assign v_STP_5101_out0 = v_EQ8_1194_out0;
assign v_JEQ_5167_out0 = v_EQ7_1608_out0;
assign v_R2_5194_out0 = v_R2_5364_out0;
assign v__5310_out0 = v_IR_1413_out0[11:10];
assign v_EXEC2LS_5403_out0 = v_EXEC2LS_1554_out0;
assign v_G1_5491_out0 = v_EQ1_156_out0 || v_EQ9_1165_out0;
assign v_4BITCOUNTERTRANSIMITER_5539_out0 = v_4BITCOUNTER_4_out0;
assign v_START_6598_out0 = v_START_1476_out0;
assign v_NORMAL_6615_out0 = v_NORMAL_93_out0;
assign v_IR_6640_out0 = v_IR_1413_out0;
assign v_9_6712_out0 = v_9_834_out0;
assign v_9_6713_out0 = v_9_835_out0;
assign v_STP_28_out0 = v_STP_5101_out0;
assign v_IR_54_out0 = v_IR_6640_out0;
assign v_G9_111_out0 = v_G6_2214_out0 || v_G7_586_out0;
assign v_START_191_out0 = v_START_6598_out0;
assign v_9_203_out0 = v_9_6713_out0;
assign v_OP_301_out0 = v__2_out0;
assign v_G7_826_out0 = v_G1_573_out0 && v_Q1_152_out0;
assign v_UART_890_out0 = v_G2_1293_out0;
assign v_G3_953_out0 = v_EQ11_1196_out0 || v_G1_5491_out0;
assign v_D_1027_out0 = v__5310_out0;
assign v_JEQ_1089_out0 = v_JEQ_5167_out0;
assign v_UARTCOUNTER_1137_out0 = v_4BITCOUNTER_1419_out0;
assign v__1181_out0 = v_IR_6640_out0[8:8];
assign v_IR15_1201_out0 = v__3482_out0;
assign v_G1_1320_out0 = v_RESET_5501_out0 && v_D_3775_out0;
assign v_G1_1324_out0 = v_RESET_5505_out0 && v_D_3779_out0;
assign v__1353_out0 = { v__1444_out0,v_Q3_5177_out0 };
assign v__1354_out0 = { v__1445_out0,v_Q3_5178_out0 };
assign v__1390_out0 = v_IR_6640_out0[4:0];
assign v_G2_1569_out0 = ! v_9_6712_out0;
assign v_EXEC2LS_1573_out0 = v_EXEC2LS_5403_out0;
assign v_JMP_1574_out0 = v_JMP_4342_out0;
assign v__1922_out0 = v_IR_6640_out0[7:4];
assign v__2361_out0 = v_IR_6640_out0[9:9];
assign v_SEL1_2842_out0 = v_IR_6640_out0[15:12];
assign v_BIT_3396_out0 = v_MUX1_314_out0;
assign v_JUMPADRESS_3419_out0 = v_ADRESS_1141_out0;
assign v_EXEC1_3451_out0 = v_EXEC1LS_3338_out0;
assign v_M_3522_out0 = v__1267_out0;
assign v_FLOAT_3772_out0 = v_FLOAT_2247_out0;
assign v_NORMAL_5057_out0 = v_NORMAL_6615_out0;
assign v_EXEC1LS_5171_out0 = v_EXEC1LS_3338_out0;
assign v_G5_5369_out0 = v_Q0_303_out0 && v_G2_3336_out0;
assign v__5494_out0 = v_IR_6640_out0[3:2];
assign v_JMI_6575_out0 = v_JMI_948_out0;
assign v_G3_6720_out0 = v_G1_573_out0 && v_G2_3336_out0;
assign v_RECEIVER_1BIT_42_out0 = v_BIT_3396_out0;
assign v_JMI_47_out0 = v_JMI_6575_out0;
assign v_B_136_out0 = v__1922_out0;
assign v_G1_138_out0 = v_EQ2_4827_out0 && v_G2_1569_out0;
assign v_STALL_208_out0 = v_G3_953_out0;
assign v__261_out0 = { v_G1_5318_out0,v_G9_111_out0 };
assign v_JMP_268_out0 = v_JMP_1574_out0;
assign v_EQ1_907_out0 = v_SEL1_2842_out0 == 4'h1;
assign v_G8_1289_out0 = ! v_9_203_out0;
assign v_EXEC2LS_1389_out0 = v_EXEC2LS_1573_out0;
assign v_G6_1415_out0 = v_G3_6720_out0 || v_G7_826_out0;
assign v_G3_1435_out0 = v_FLOAT_3772_out0 && v_NORMAL_6615_out0;
assign v_EQ3_1447_out0 = v_SEL1_2842_out0 == 4'h9;
assign v_EXEC2_1545_out0 = v_NORMAL_5057_out0;
assign v_JMI_1565_out0 = v_JMI_6575_out0;
assign v_JEQ_2174_out0 = v_JEQ_1089_out0;
assign v_JUMPADRESS_2316_out0 = v_JUMPADRESS_3419_out0;
assign v_K_2838_out0 = v__1390_out0;
assign v_JMP_3475_out0 = v_JMP_1574_out0;
assign v_C_4259_out0 = v__2361_out0;
assign v_SHIFT_4263_out0 = v__5494_out0;
assign v_D_4307_out0 = v_D_1027_out0;
assign v_JEQ_4334_out0 = v_JEQ_1089_out0;
assign v_STP_5154_out0 = v_STP_28_out0;
assign v_AD2_5266_out0 = v_M_3522_out0;
assign v_EXEC1_5298_out0 = v_EXEC1_3451_out0;
assign v_IR_5321_out0 = v_IR_54_out0;
assign v_UART_5325_out0 = v_UART_890_out0;
assign v_UART_COUNTER_5328_out0 = v_UARTCOUNTER_1137_out0;
assign v_EXEC1LS_5335_out0 = v_EXEC1LS_5171_out0;
assign v_STP_5402_out0 = v_STP_28_out0;
assign v_OP_5524_out0 = v_OP_301_out0;
assign v_S_5562_out0 = v__1181_out0;
assign v_8BITCOUNTER_6549_out0 = v__1353_out0;
assign v_8BITCOUNTER_6550_out0 = v__1354_out0;
assign v_EQ2_6752_out0 = v_SEL1_2842_out0 == 4'h2;
assign v_AD1_6785_out0 = v_D_1027_out0;
assign v_B_567_out0 = v_B_136_out0;
assign v_EQ6_827_out0 = v_OP_5524_out0 == 3'h5;
assign v__845_out0 = v_IR_5321_out0[14:14];
assign v_STALL_860_out0 = v_STALL_208_out0;
assign v_G15_906_out0 = !(v_EXEC1_5298_out0 || v_FF1_26_out0);
assign v_EXEC2_982_out0 = v_EXEC2_1545_out0;
assign v_RD_1006_out0 = v_D_4307_out0;
assign v_EQ4_1047_out0 = v_8BITCOUNTER_6549_out0 == 4'h0;
assign v__1185_out0 = v_IR_5321_out0[15:15];
assign v_IN_1202_out0 = v_RECEIVER_1BIT_42_out0;
assign v__1204_out0 = v_IR_5321_out0[13:13];
assign v_K_1285_out0 = v_K_2838_out0;
assign v_EXEC2_1290_out0 = v_EXEC2LS_1389_out0;
assign v_JMP_1301_out0 = v_JMP_3475_out0;
assign v_SUB_1315_out0 = v_EQ3_1447_out0;
assign v__1382_out0 = v_AD2_5266_out0[0:0];
assign v__1382_out1 = v_AD2_5266_out0[1:1];
assign v__1396_out0 = v_IR_5321_out0[12:12];
assign v_EQ8_1440_out0 = v_OP_5524_out0 == 3'h7;
assign v_MULTI_OPCODE_1474_out0 = v_EQ1_907_out0;
assign v_EXEC2LS_1503_out0 = v_EXEC2LS_1389_out0;
assign v__1899_out0 = v_IR_5321_out0[9:0];
assign v__1899_out1 = v_IR_5321_out0[15:6];
assign v_G3_1932_out0 = v_EQ2_6752_out0 && v_FLOATING_INS_6796_out0;
assign v_EXEC1LS_2293_out0 = v_EXEC1LS_5335_out0;
assign v__3376_out0 = v_AD1_6785_out0[0:0];
assign v__3376_out1 = v_AD1_6785_out0[1:1];
assign v_STALL_3392_out0 = v_STALL_208_out0;
assign v_EQ1_3483_out0 = v_OP_5524_out0 == 3'h0;
assign v_EQ3_3495_out0 = v_OP_5524_out0 == 3'h2;
assign v_EXEC1_3496_out0 = v_EXEC1LS_5335_out0;
assign v_JMI_4273_out0 = v_JMI_47_out0;
assign v_EQ1_5091_out0 = v_8BITCOUNTER_6550_out0 == 4'h0;
assign v_EQ4_5098_out0 = v_OP_5524_out0 == 3'h3;
assign v_EQ5_5106_out0 = v_OP_5524_out0 == 3'h4;
assign v_EQ7_5122_out0 = v_OP_5524_out0 == 3'h6;
assign v_UART_5176_out0 = v_UART_5325_out0;
assign v_SHIFT_5225_out0 = v_SHIFT_4263_out0;
assign v_EQ2_5301_out0 = v_OP_5524_out0 == 3'h1;
assign v_8BITCOUNTER_5462_out0 = v_8BITCOUNTER_6549_out0;
assign v_STP_5531_out0 = v_STP_5154_out0;
assign v_STP_6646_out0 = v_STP_5402_out0;
assign v_JEQ_6682_out0 = v_JEQ_2174_out0;
assign v_C_6782_out0 = v_C_4259_out0;
assign v_BIT_STREAM_IN_7_out0 = v_IN_1202_out0;
assign v__64_out0 = { v_K_1285_out0,v_C1_294_out0 };
assign v_G5_102_out0 = !(v_EQ2_5404_out0 && v_EQ1_5091_out0);
assign v_C_118_out0 = v_C_6782_out0;
assign v_MUX4_186_out0 = v__1382_out0 ? v_R1_4311_out0 : v_R0_828_out0;
assign v_EXEC2_215_out0 = v_EXEC2_982_out0;
assign v_FLOATING_EN_ALU_307_out0 = v_G3_1932_out0;
assign v_G9_821_out0 = ! v_STALL_3392_out0;
assign v_EXEC1_910_out0 = v_EXEC1LS_2293_out0;
assign v_MUX1_1235_out0 = v__3376_out0 ? v_REG1_1128_out0 : v_REG0_5368_out0;
assign v_NOTUSED_1317_out0 = v__1899_out1;
assign v_SUB_INSTRUCTION_1361_out0 = v_SUB_1315_out0;
assign v_EXEC1_1481_out0 = v_EXEC1_3496_out0;
assign v_EXEC2_1578_out0 = v_EXEC2LS_1503_out0;
assign v_TST_1861_out0 = v_EQ8_1440_out0;
assign v_AND_1880_out0 = v_EQ7_5122_out0;
assign v_UART_1897_out0 = v_UART_5176_out0;
assign v_MULTI_INSTRUCTION_1928_out0 = v_MULTI_OPCODE_1474_out0;
assign v_G24_1930_out0 = ! v__1204_out0;
assign v_ADD_2179_out0 = v_EQ1_3483_out0;
assign v__2211_out0 = v__1899_out0[8:0];
assign v__2211_out1 = v__1899_out0[9:1];
assign v_MUX2_2252_out0 = v__3376_out0 ? v_REG3_2317_out0 : v_REG2_6035_out0;
assign v_BIN_2868_out0 = v_B_567_out0;
assign v_G28_3373_out0 = ! v__845_out0;
assign v_G25_3418_out0 = v__1185_out0 && v__845_out0;
assign v_G6_3443_out0 = !(v_EQ5_4313_out0 && v_EQ4_1047_out0);
assign v_EXEC2_3524_out0 = v_EXEC2_1290_out0;
assign v_SUB_4264_out0 = v_EQ2_5301_out0;
assign v_MUX5_4349_out0 = v__1382_out0 ? v_R3_2273_out0 : v_R2_1484_out0;
assign v_STALL_5070_out0 = v_STALL_860_out0;
assign v_G4_5071_out0 = v_G5_5369_out0 && v_STALL_3392_out0;
assign v_MOV_5117_out0 = v_EQ5_5106_out0;
assign v_ADC_5119_out0 = v_EQ3_3495_out0;
assign v_G12_5202_out0 = ! v_STP_5531_out0;
assign v_EXEC1LS_5268_out0 = v_EXEC1LS_2293_out0;
assign v_G5_5408_out0 = ! v_EQ4_1047_out0;
assign v_MULTI_OPCODE_5461_out0 = v_MULTI_OPCODE_1474_out0;
assign v_G6_5508_out0 = ! v_EQ1_5091_out0;
assign v_G2_6027_out0 = v_EXEC2_982_out0 || v_EXEC2LS_1503_out0;
assign v_G11_6620_out0 = v_EXEC1_5298_out0 || v_STP_5531_out0;
assign v_G9_6684_out0 = v_EQ2_5404_out0 && v_EQ1_5091_out0;
assign v_SBC_6705_out0 = v_EQ4_5098_out0;
assign v_CMP_6707_out0 = v_EQ6_827_out0;
assign v_G8_9_out0 = v_G1_138_out0 && v_BIT_STREAM_IN_7_out0;
assign v_EXEC1_12_out0 = v_EXEC1_910_out0;
assign v_MOV_99_out0 = v_MOV_5117_out0;
assign v_MUX3_155_out0 = v__3376_out1 ? v_MUX2_2252_out0 : v_MUX1_1235_out0;
assign v_C_187_out0 = v_C_118_out0;
assign v_MUX1_262_out0 = v_C_118_out0 ? v_ROR_34_out0 : v_SHIFT_5225_out0;
assign v_MUX2_562_out0 = v_G2_6027_out0 ? v_D_1027_out0 : v_M_3522_out0;
assign v_EQ1_568_out0 = v__2211_out1 == 1'h0;
assign v_TRANSMITER_OVERFLOW_830_out0 = v_G6_5508_out0;
assign v_OVERFLOW_RX_858_out0 = v_G6_3443_out0;
assign v_G8_863_out0 = v_G7_826_out0 || v_G4_5071_out0;
assign v_TX_IN_PROGRESS_911_out0 = v_G5_102_out0;
assign v_G1_1085_out0 = ! v_TST_1861_out0;
assign v_BIT_1135_out0 = v_BIT_STREAM_IN_7_out0;
assign v_MUX6_1142_out0 = v__1382_out1 ? v_MUX5_4349_out0 : v_MUX4_186_out0;
assign v_G7_1195_out0 = v_G9_6684_out0 || v_G8_1289_out0;
assign v_G11_1280_out0 = v_G5_5369_out0 && v_G9_821_out0;
assign v_EXEC1_1284_out0 = v_EXEC1LS_5268_out0;
assign v_G23_1387_out0 = v_G25_3418_out0 && v_G24_1930_out0;
assign v_SUB_1417_out0 = v_G11_6620_out0;
assign v_SUB_1442_out0 = v_SUB_4264_out0;
assign v_CMP_1855_out0 = v_CMP_6707_out0;
assign v_SBC_2356_out0 = v_SBC_6705_out0;
assign v_G2_3380_out0 = v_S_5562_out0 && v_EXEC2_215_out0;
assign v_STARTBIT_3420_out0 = v_BIT_STREAM_IN_7_out0;
assign v_EQ2_3481_out0 = v__2211_out1 == 1'h1;
assign v_MULTI_OPCODE_3499_out0 = v_MULTI_OPCODE_5461_out0;
assign v_TST_4300_out0 = v_TST_1861_out0;
assign v_G27_4825_out0 = v__1185_out0 && v_G28_3373_out0;
assign v_G5_5142_out0 = ! v_CMP_6707_out0;
assign v_G3_5151_out0 = v_EQ6_11_out0 && v_G5_5408_out0;
assign v__5347_out0 = v__2211_out0[7:0];
assign v__5347_out1 = v__2211_out0[8:1];
assign v_uart_5478_out0 = v_UART_1897_out0;
assign v_ADD_5509_out0 = v_ADD_2179_out0;
assign v_SUB_INSTRUCTION_5510_out0 = v_SUB_INSTRUCTION_1361_out0;
assign v__6536_out0 = v_BIN_2868_out0[3:1];
assign v_MULTI_INSTRUCTION_6565_out0 = v_MULTI_INSTRUCTION_1928_out0;
assign v_KEXTEND_6567_out0 = v__64_out0;
assign v_AND_6681_out0 = v_AND_1880_out0;
assign v_ADC_6710_out0 = v_ADC_5119_out0;
assign v_G3_10_out0 = v_G1_1085_out0 && v_EXEC2_215_out0;
assign v_RX_OVERFLOW_15_out0 = v_OVERFLOW_RX_858_out0;
assign v_G5_114_out0 = ((v__1590_out0 && !v_SUB_1417_out0) || (!v__1590_out0) && v_SUB_1417_out0);
assign v_SR_184_out0 = v_MUX1_262_out0;
assign v_TST_198_out0 = v_TST_4300_out0;
assign v_SR_266_out0 = v_MUX1_262_out0;
assign v_MULTI_INSTRUCTION_300_out0 = v_MULTI_INSTRUCTION_6565_out0;
assign v_STORE_585_out0 = v_EQ1_568_out0;
assign v_DOUT1_591_out0 = v_MUX3_155_out0;
assign v_DOUT2_848_out0 = v_MUX6_1142_out0;
assign v_ADC_889_out0 = v_ADC_6710_out0;
assign v_SR_957_out0 = v_MUX1_262_out0;
assign v_G8_987_out0 = ((v__88_out0 && !v_SUB_1417_out0) || (!v__88_out0) && v_SUB_1417_out0);
assign v__1045_out0 = { v_C1_5309_out0,v__6536_out0 };
assign v_G9_1138_out0 = ((v__1106_out0 && !v_SUB_1417_out0) || (!v__1106_out0) && v_SUB_1417_out0);
assign v_G6_1178_out0 = ((v__986_out0 && !v_SUB_1417_out0) || (!v__986_out0) && v_SUB_1417_out0);
assign v_MULTI_INSTRUCTION_1193_out0 = v_MULTI_INSTRUCTION_6565_out0;
assign v_G11_1243_out0 = ((v__31_out0 && !v_SUB_1417_out0) || (!v__31_out0) && v_SUB_1417_out0);
assign v_G3_1277_out0 = ((v__142_out0 && !v_SUB_1417_out0) || (!v__142_out0) && v_SUB_1417_out0);
assign v_G10_1283_out0 = ((v__5532_out0 && !v_SUB_1417_out0) || (!v__5532_out0) && v_SUB_1417_out0);
assign v_tx_Overflow_1349_out0 = v_TRANSMITER_OVERFLOW_830_out0;
assign v_G2_1408_out0 = v_EXEC1_1284_out0 && v_G3_843_out0;
assign v_tx_in_progress_1449_out0 = v_TX_IN_PROGRESS_911_out0;
assign v__1482_out0 = { v__1443_out1,v_BIT_1135_out0 };
assign v_LOAD_1519_out0 = v_EQ2_3481_out0;
assign v_G2_1577_out0 = ((v__1523_out0 && !v_SUB_1417_out0) || (!v__1523_out0) && v_SUB_1417_out0);
assign v_G12_2294_out0 = ((v__917_out0 && !v_SUB_1417_out0) || (!v__917_out0) && v_SUB_1417_out0);
assign v_G26_2312_out0 = v_G23_1387_out0 && v__1396_out0;
assign v_G7_2354_out0 = ((v__6599_out0 && !v_SUB_1417_out0) || (!v__6599_out0) && v_SUB_1417_out0);
assign v_W_EN_3377_out0 = v__5347_out1;
assign v__3467_out0 = v__5347_out0[6:0];
assign v__3467_out1 = v__5347_out0[7:1];
assign v_SUB_INSTRUCTION_3478_out0 = v_SUB_INSTRUCTION_5510_out0;
assign v_CMP_4255_out0 = v_CMP_1855_out0;
assign v_G12_5088_out0 = v_G11_1280_out0 && v_G2_3336_out0;
assign v_G7_5093_out0 = v_9_6712_out0 && v_G3_5151_out0;
assign v_G35_5104_out0 = v_STARTBIT_3420_out0 && v_G36_1528_out0;
assign v_G1_5159_out0 = ((v__6683_out0 && !v_SUB_1417_out0) || (!v__6683_out0) && v_SUB_1417_out0);
assign v_AD3_5161_out0 = v_MUX2_562_out0;
assign v_SR_5221_out0 = v_MUX1_262_out0;
assign v_SBC_5438_out0 = v_SBC_2356_out0;
assign v_BYTERECEIVED_5511_out0 = v_G8_9_out0;
assign v_G4_6030_out0 = ((v__92_out0 && !v_SUB_1417_out0) || (!v__92_out0) && v_SUB_1417_out0);
assign v_SUB_6033_out0 = v_SUB_1442_out0;
assign v_AD3_6545_out0 = v_MUX2_562_out0;
assign v_LOAD_115_out0 = v_LOAD_1519_out0;
assign v_ROR_140_out0 = v_SR_266_out0 == 2'h3;
assign v_G6_162_out0 = v_C_1559_out0 && v_ADC_889_out0;
assign v_G9_197_out0 = ! v_W_EN_3377_out0;
assign v_G9_199_out0 = ((v_AND_6681_out0 && !v_TST_198_out0) || (!v_AND_6681_out0) && v_TST_198_out0);
assign v_LSR_204_out0 = v_SR_184_out0 == 2'h1;
assign v_G5_221_out0 = v_STORE_585_out0 && v_EXEC1_12_out0;
assign v_RD_245_out0 = v_DOUT1_591_out0;
assign v_STORE_265_out0 = v_STORE_585_out0;
assign v_ROR_267_out0 = v_SR_184_out0 == 2'h3;
assign v_LSR_576_out0 = v_SR_266_out0 == 2'h1;
assign v__836_out0 = { v_G1_5159_out0,v_G2_1577_out0 };
assign v_G10_857_out0 = v_G6_1415_out0 || v_G12_5088_out0;
assign v_ENABLE_859_out0 = v_G7_5093_out0;
assign v_LSL_909_out0 = v_SR_266_out0 == 2'h0;
assign v_G2_923_out0 = v_W_EN_3377_out0 && v_EXEC1_12_out0;
assign v_ENABLE_984_out0 = v_G35_5104_out0;
assign v_MUX1_1174_out0 = v_C_187_out0 ? v__1045_out0 : v_BIN_2868_out0;
assign v_LSL_1388_out0 = v_SR_5221_out0 == 2'h0;
assign v_G3_1414_out0 = v_LOAD_1519_out0 && v_EXEC2_3524_out0;
assign v_G1_1473_out0 = v_SBC_5438_out0 && v_C_1559_out0;
assign v_LSL_1486_out0 = v_SR_184_out0 == 2'h0;
assign v_LSL_1551_out0 = v_SR_957_out0 == 2'h0;
assign v_ROR_1598_out0 = v_SR_5221_out0 == 2'h3;
assign v_ROR_1599_out0 = v_SR_957_out0 == 2'h3;
assign v_TX_OVERFLOW_1902_out0 = v_tx_Overflow_1349_out0;
assign v_tx_in_progress_1925_out0 = v_tx_in_progress_1449_out0;
assign v_G5_2187_out0 = v_SUB_6033_out0 || v_CMP_4255_out0;
assign v_G4_2313_out0 = ((v_SBC_5438_out0 && !v_ADC_889_out0) || (!v_SBC_5438_out0) && v_ADC_889_out0);
assign v_G29_2860_out0 = v_G26_2312_out0 || v_G27_4825_out0;
assign v_LSR_3393_out0 = v_SR_957_out0 == 2'h1;
assign v_G3_4265_out0 = ((v_SUB_6033_out0 && !v_CMP_4255_out0) || (!v_SUB_6033_out0) && v_CMP_4255_out0);
assign v_AD3_4269_out0 = v_AD3_6545_out0;
assign v_ASR_4308_out0 = v_SR_957_out0 == 2'h2;
assign v_ASR_5107_out0 = v_SR_266_out0 == 2'h2;
assign v__5164_out0 = v__3467_out0[5:0];
assign v__5164_out1 = v__3467_out0[6:1];
assign v_ASR_5199_out0 = v_SR_184_out0 == 2'h2;
assign v_done_receiving_5219_out0 = v_BYTERECEIVED_5511_out0;
assign v_P_5258_out0 = v__3467_out1;
assign v_RX_OVERFLOW_5535_out0 = v_RX_OVERFLOW_15_out0;
assign v_G4_6032_out0 = v_G5_5142_out0 && v_G3_10_out0;
assign v_MULTI_INSTRUCTION_6558_out0 = v_MULTI_INSTRUCTION_300_out0;
assign v_LSR_6568_out0 = v_SR_5221_out0 == 2'h1;
assign v_RM_6701_out0 = v_DOUT2_848_out0;
assign v_ASR_6755_out0 = v_SR_5221_out0 == 2'h2;
assign v_RM_6773_out0 = v_DOUT2_848_out0;
assign v_G1_6786_out0 = v_G2_1408_out0 || v_EXEC2_1578_out0;
assign v_G4_109_out0 = v_G2_923_out0 || v_G3_1414_out0;
assign v__559_out0 = v__5164_out0[1:0];
assign v__559_out1 = v__5164_out0[5:4];
assign v_G1_583_out0 = ! v__5164_out1;
assign v__1163_out0 = { v__836_out0,v_G3_1277_out0 };
assign v_RDOUT_1360_out0 = v_RD_245_out0;
assign v_LOAD_1412_out0 = v_LOAD_115_out0;
assign v_RD_1896_out0 = v_RD_245_out0;
assign v_OP1_1900_out0 = v_RD_245_out0;
assign v_G8_2178_out0 = v_G1_1473_out0 || v_G6_162_out0;
assign v_G7_2186_out0 = v_P_5258_out0 && v_EXEC1_12_out0;
assign v_G10_2188_out0 = v_EXEC2_3524_out0 && v_P_5258_out0;
assign v_RM_2217_out0 = v_RM_6773_out0;
assign v_EN_2243_out0 = v_G29_2860_out0;
assign v_DONE_RECEIVING_3470_out0 = v_done_receiving_5219_out0;
assign v_G5_3486_out0 = v_MULTI_INSTRUCTION_6558_out0 || v_DIV_INSTRUCTION_2254_out0;
assign v_RM_4298_out0 = v_RM_6773_out0;
assign v_G18_4330_out0 = !(v_ENABLE_984_out0 || v_Q7_3382_out0);
assign v_MUX1_4337_out0 = v_C_4259_out0 ? v_KEXTEND_6567_out0 : v_RM_6701_out0;
assign v_TX_IN_PROG_5059_out0 = v_tx_in_progress_1925_out0;
assign v_MUX10_5120_out0 = v_MULTI_INSTRUCTION_6558_out0 ? v_C13_196_out0 : v_C12_1029_out0;
assign v_RAMWEN_5267_out0 = v_G5_221_out0;
assign v_B_5311_out0 = v_MUX1_1174_out0;
assign v_STORE_5329_out0 = v_STORE_265_out0;
assign v_WENALU_5345_out0 = v_G4_6032_out0;
assign v_G2_5481_out0 = ((v_ADD_5509_out0 && !v_G3_4265_out0) || (!v_ADD_5509_out0) && v_G3_4265_out0);
assign v_G11_5495_out0 = v_G5_2187_out0 || v_SBC_5438_out0;
assign v_RM_5496_out0 = v_RM_6773_out0;
assign v_WENMULTI_5515_out0 = v_G1_6786_out0;
assign v_G14_6542_out0 = v_G10_857_out0 || v_G13_3477_out0;
assign v_G4_6750_out0 = ! v_MULTI_INSTRUCTION_6558_out0;
assign v_SEL6_53_out0 = v_RM_5496_out0[9:0];
assign v_G10_67_out0 = v_G8_2178_out0 || v_G5_2187_out0;
assign v_G7_87_out0 = ((v_G2_5481_out0 && !v_G4_2313_out0) || (!v_G2_5481_out0) && v_G4_2313_out0);
assign v__94_out0 = v_B_5311_out0[3:3];
assign v__201_out0 = v_B_5311_out0[1:1];
assign v__846_out0 = v_B_5311_out0[0:0];
assign v_G9_1046_out0 = v_DONE_RECEIVING_3470_out0 && v_Q_3786_out0;
assign v_WENRAM_1134_out0 = v_RAMWEN_5267_out0;
assign v_WEN_MULTI_1164_out0 = v_WENMULTI_5515_out0;
assign v_SEL3_1274_out0 = v_RD_1896_out0[15:15];
assign v_G8_1278_out0 = v_G9_197_out0 && v_G10_2188_out0;
assign v_SEL1_1421_out0 = v_RD_1896_out0[14:10];
assign v__1448_out0 = { v__1163_out0,v_G4_6030_out0 };
assign v_OP1_1454_out0 = v_OP1_1900_out0;
assign v_RM_1555_out0 = v_RM_4298_out0;
assign v_G21_1856_out0 = v_G18_4330_out0 || v_G22_5405_out0;
assign v_SUB_2255_out0 = v_G11_5495_out0;
assign v_M_2295_out0 = v__559_out0;
assign v_LOAD_3488_out0 = v_LOAD_1412_out0;
assign v_SEL4_3752_out0 = v_RM_5496_out0[15:15];
assign v_N_3755_out0 = v__559_out1;
assign v_WENALU_4262_out0 = v_WENALU_5345_out0;
assign v_SEL5_4314_out0 = v_RD_1896_out0[9:0];
assign v_BYTE_READY_RX_4826_out0 = v_DONE_RECEIVING_3470_out0;
assign v_REGISTER_OUT_5064_out0 = v_RDOUT_1360_out0;
assign v_U_5155_out0 = v_G1_583_out0;
assign v__5308_out0 = v_B_5311_out0[2:2];
assign v__5441_out0 = { v_G14_6542_out0,v_G8_863_out0 };
assign v_IN_5542_out0 = v_MUX1_4337_out0;
assign v_STORE_6555_out0 = v_STORE_5329_out0;
assign v_SEL2_6566_out0 = v_RM_5496_out0[14:10];
assign v_G6_6648_out0 = v_DONE_RECEIVING_3470_out0 || v_Q_3786_out0;
assign v_RM_6657_out0 = v_RM_2217_out0;
assign v_WENLDST_6775_out0 = v_G4_109_out0;
assign v_IN_51_out0 = v_IN_5542_out0;
assign v_STORE_110_out0 = v_STORE_6555_out0;
assign v_RAM_IN_116_out0 = v_REGISTER_OUT_5064_out0;
assign v_RD_SIGN_141_out0 = v_SEL3_1274_out0;
assign v_D_302_out0 = v__5441_out0;
assign v_RD_SIG_865_out0 = v_SEL5_4314_out0;
assign v_OP1_1005_out0 = v_OP1_1454_out0;
assign v_EN_1136_out0 = v__846_out0;
assign v_EN_1190_out0 = v__94_out0;
assign v_OP2_EXP_1242_out0 = v_SEL2_6566_out0;
assign v_WENLDST_1309_out0 = v_WENLDST_6775_out0;
assign v__1479_out0 = v_RM_6657_out0[11:0];
assign v__1479_out1 = v_RM_6657_out0[15:4];
assign v_BYTE_READY_2239_out0 = v_BYTE_READY_RX_4826_out0;
assign v_SUB_2256_out0 = v_U_5155_out0;
assign v_WENRAM_2272_out0 = v_WENRAM_1134_out0;
assign v__2866_out0 = { v__1448_out0,v_G5_114_out0 };
assign v_LOAD_4312_out0 = v_LOAD_3488_out0;
assign v_RD_EXP_4352_out0 = v_SEL1_1421_out0;
assign v_WEN_MULTI_5113_out0 = v_WEN_MULTI_1164_out0;
assign v_EN_5158_out0 = v__201_out0;
assign v_OP2_SIGN_5333_out0 = v_SEL4_3752_out0;
assign v__5527_out0 = { v_N_3755_out0,v_C1_1564_out0 };
assign v_EN_6500_out0 = v__5308_out0;
assign v_G6_6537_out0 = v_G8_1278_out0 || v_G7_2186_out0;
assign v_OP2_SIG_6556_out0 = v_SEL6_53_out0;
assign v_REGISTER_OUTPUT_6728_out0 = v_REGISTER_OUT_5064_out0;
assign v__50_out0 = { v__2866_out0,v_G6_1178_out0 };
assign v_split_214_out0 = v_REGISTER_OUTPUT_6728_out0[7:0];
assign v_split_214_out1 = v_REGISTER_OUTPUT_6728_out0[15:8];
assign v_OP2_EXP_263_out0 = v_OP2_EXP_1242_out0;
assign v_SIG_RM_864_out0 = v_OP2_SIG_6556_out0;
assign v_RD_SIGN_1173_out0 = v_RD_SIGN_141_out0;
assign v_WRITE_EN_1582_out0 = v_WENRAM_2272_out0;
assign v_RD_EXP_1927_out0 = v_RD_EXP_4352_out0;
assign v_WEN_MULTI_2240_out0 = v_WEN_MULTI_5113_out0;
assign v__2248_out0 = v_D_302_out0[0:0];
assign v__2248_out1 = v_D_302_out0[1:1];
assign v_EXP_RM_2315_out0 = v_OP2_EXP_1242_out0;
assign v__2358_out0 = v_IN_51_out0[14:0];
assign v__2358_out1 = v_IN_51_out0[15:1];
assign v_EXP_RD_2869_out0 = v_RD_EXP_4352_out0;
assign v_MUX3_4339_out0 = v_IR15_1201_out0 ? v_WENALU_4262_out0 : v_WENLDST_1309_out0;
assign v_A_5067_out0 = v_OP1_1005_out0;
assign v_BYTE_READY_5498_out0 = v_BYTE_READY_2239_out0;
assign v_OP2_SIGN_5516_out0 = v_OP2_SIGN_5333_out0;
assign v_A_5538_out0 = v__5527_out0;
assign v_SIG_RD_5561_out0 = v_RD_SIG_865_out0;
assign v_UNUSED_6616_out0 = v__1479_out1;
assign v_BYTE_READY_RX_6654_out0 = v_BYTE_READY_2239_out0;
assign v_IN_6792_out0 = v_IN_51_out0;
assign v__1_out0 = v_A_5067_out0[4:4];
assign v__37_out0 = { v__50_out0,v_G7_2354_out0 };
assign v__41_out0 = v_A_5538_out0[3:3];
assign v__98_out0 = v_A_5538_out0[15:15];
assign v_G1_143_out0 = ((v_OP2_SIGN_5516_out0 && !v_SUB_INSTRUCTION_3478_out0) || (!v_OP2_SIGN_5516_out0) && v_SUB_INSTRUCTION_3478_out0);
assign v__160_out0 = v_A_5538_out0[0:0];
assign v__164_out0 = v_A_5538_out0[9:9];
assign v__832_out0 = v_A_5067_out0[5:5];
assign v__854_out0 = v_A_5067_out0[11:11];
assign v__927_out0 = v_A_5067_out0[0:0];
assign v__1023_out0 = v_A_5538_out0[13:13];
assign v__1049_out0 = v_A_5067_out0[2:2];
assign v__1180_out0 = v_A_5538_out0[6:6];
assign v_RD_EXP_1268_out0 = v_RD_EXP_1927_out0;
assign v__1348_out0 = v_A_5067_out0[15:15];
assign v__1402_out0 = v_A_5067_out0[12:12];
assign v__1404_out0 = v_A_5067_out0[3:3];
assign v__1522_out0 = v_A_5538_out0[14:14];
assign v__1581_out0 = v_A_5067_out0[8:8];
assign v__1597_out0 = v_A_5538_out0[2:2];
assign v__2245_out0 = v_A_5067_out0[10:10];
assign v__2301_out0 = v_A_5067_out0[13:13];
assign v_BYTE_READY_3447_out0 = v_BYTE_READY_5498_out0;
assign v__3523_out0 = { v_C1_293_out0,v__2358_out0 };
assign v__4306_out0 = v_A_5538_out0[8:8];
assign v_MUX6_4309_out0 = v_MULTI_OPCODE_1474_out0 ? v_WEN_MULTI_1164_out0 : v_MUX3_4339_out0;
assign v__4344_out0 = v_A_5538_out0[7:7];
assign v__4354_out0 = v_A_5067_out0[14:14];
assign v_EQ2_5099_out0 = v_EXP_RM_2315_out0 == 5'h0;
assign v__5112_out0 = v_A_5538_out0[5:5];
assign v_OP2_EXP_5114_out0 = v_OP2_EXP_263_out0;
assign v__5116_out0 = v_A_5538_out0[1:1];
assign v__5265_out0 = v_A_5538_out0[4:4];
assign v__5305_out0 = v_A_5538_out0[12:12];
assign v__5344_out0 = v_A_5538_out0[10:10];
assign v__5488_out0 = v_A_5067_out0[6:6];
assign v_UNNOTUSED_5522_out0 = v__2358_out1;
assign v__6594_out0 = v_A_5067_out0[7:7];
assign v_EQ1_6617_out0 = v_EXP_RD_2869_out0 == 5'h0;
assign v__6660_out0 = v_A_5067_out0[1:1];
assign v__6680_out0 = v_A_5538_out0[11:11];
assign v__6715_out0 = v_A_5067_out0[9:9];
assign v_MUX1_19_out0 = v_LSL_1551_out0 ? v__3523_out0 : v_IN_6792_out0;
assign v_G3_104_out0 = ((v__1597_out0 && !v_SUB_2256_out0) || (!v__1597_out0) && v_SUB_2256_out0);
assign v_G1_312_out0 = ! v_EQ1_6617_out0;
assign v_G8_596_out0 = ((v__4344_out0 && !v_SUB_2256_out0) || (!v__4344_out0) && v_SUB_2256_out0);
assign v_WEN3_829_out0 = v_MUX6_4309_out0;
assign v_EQ2_856_out0 = v_OP2_EXP_5114_out0 == 5'h0;
assign v_G15_887_out0 = ((v__1522_out0 && !v_SUB_2256_out0) || (!v__1522_out0) && v_SUB_2256_out0);
assign v_EQ1_1266_out0 = v_RD_EXP_1268_out0 == 5'h0;
assign v_G7_1357_out0 = ((v__1180_out0 && !v_SUB_2256_out0) || (!v__1180_out0) && v_SUB_2256_out0);
assign v_G12_1627_out0 = ((v__6680_out0 && !v_SUB_2256_out0) || (!v__6680_out0) && v_SUB_2256_out0);
assign v_G14_2216_out0 = ((v__1023_out0 && !v_SUB_2256_out0) || (!v__1023_out0) && v_SUB_2256_out0);
assign v_G13_2298_out0 = ((v__5305_out0 && !v_SUB_2256_out0) || (!v__5305_out0) && v_SUB_2256_out0);
assign v_G2_3444_out0 = ! v_EQ2_5099_out0;
assign v_G2_3450_out0 = ((v__5116_out0 && !v_SUB_2256_out0) || (!v__5116_out0) && v_SUB_2256_out0);
assign v__4274_out0 = { v__37_out0,v_G8_987_out0 };
assign v_BYTE_READY_5195_out0 = v_BYTE_READY_3447_out0;
assign v_G5_5201_out0 = ((v__5265_out0 && !v_SUB_2256_out0) || (!v__5265_out0) && v_SUB_2256_out0);
assign v_G1_5271_out0 = v_WRITE_EN_1582_out0 || v_BYTE_READY_3447_out0;
assign v_G4_5413_out0 = ((v__41_out0 && !v_SUB_2256_out0) || (!v__41_out0) && v_SUB_2256_out0);
assign v_G16_5431_out0 = ((v__98_out0 && !v_SUB_2256_out0) || (!v__98_out0) && v_SUB_2256_out0);
assign v_G10_6518_out0 = ((v__164_out0 && !v_SUB_2256_out0) || (!v__164_out0) && v_SUB_2256_out0);
assign v_G9_6552_out0 = ((v__4306_out0 && !v_SUB_2256_out0) || (!v__4306_out0) && v_SUB_2256_out0);
assign v_G11_6573_out0 = ((v__5344_out0 && !v_SUB_2256_out0) || (!v__5344_out0) && v_SUB_2256_out0);
assign v_G6_6719_out0 = ((v__5112_out0 && !v_SUB_2256_out0) || (!v__5112_out0) && v_SUB_2256_out0);
assign v_G1_6777_out0 = ((v__160_out0 && !v_SUB_2256_out0) || (!v__160_out0) && v_SUB_2256_out0);
assign v__955_out0 = { v_G1_6777_out0,v_G2_3450_out0 };
assign v__1352_out0 = { v_SIG_RM_864_out0,v_G2_3444_out0 };
assign v__1386_out0 = { v__4274_out0,v_G9_1138_out0 };
assign v_BYTE_READY_1393_out0 = v_BYTE_READY_5195_out0;
assign v__2370_out0 = v_MUX1_19_out0[0:0];
assign v__2370_out1 = v_MUX1_19_out0[15:15];
assign v__3790_out0 = { v_SIG_RD_5561_out0,v_G1_312_out0 };
assign v_D1_4350_out0 = (v_AD3_5161_out0 == 2'b00) ? v_WEN3_829_out0 : 1'h0;
assign v_D1_4350_out1 = (v_AD3_5161_out0 == 2'b01) ? v_WEN3_829_out0 : 1'h0;
assign v_D1_4350_out2 = (v_AD3_5161_out0 == 2'b10) ? v_WEN3_829_out0 : 1'h0;
assign v_D1_4350_out3 = (v_AD3_5161_out0 == 2'b11) ? v_WEN3_829_out0 : 1'h0;
assign v_MUX13_6724_out0 = v_EQ1_1266_out0 ? v_0B00001_5193_out0 : v_RD_EXP_1268_out0;
assign v_MUX12_6789_out0 = v_EQ2_856_out0 ? v_0B00001_5193_out0 : v_OP2_EXP_5114_out0;
assign v_NOTUSED_962_out0 = v__2370_out0;
assign v__1291_out0 = { v__1386_out0,v_G10_1283_out0 };
assign v_SIG_RD_11bit_1605_out0 = v__3790_out0;
assign v_SIG_RM_11bit_3384_out0 = v__1352_out0;
assign v__4832_out0 = { v__955_out0,v_G3_104_out0 };
assign v__5061_out0 = { v_MUX13_6724_out0,v_0_5269_out0 };
assign v__5320_out0 = { v__2370_out1,v_C1_293_out0 };
assign v__5341_out0 = { v_MUX12_6789_out0,v_0_5269_out0 };
assign v_OP2_SIG11_8_out0 = v_SIG_RM_11bit_3384_out0;
assign v_XOR3_1241_out0 = v_NEG1_3398_out0 ^ v__5341_out0;
assign v_MUX2_1585_out0 = v_LSR_3393_out0 ? v__5320_out0 : v_MUX1_19_out0;
assign v__2311_out0 = { v__1291_out0,v_G11_1243_out0 };
assign v__4277_out0 = { v__4832_out0,v_G4_5413_out0 };
assign v_RD_SIG11_4356_out0 = v_SIG_RD_11bit_1605_out0;
assign v__1584_out0 = { v__4277_out0,v_G5_5201_out0 };
assign v_MUX8_2238_out0 = v_MULTI_INSTRUCTION_6558_out0 ? v__5341_out0 : v_XOR3_1241_out0;
assign v_OP2_SIG11_2357_out0 = v_OP2_SIG11_8_out0;
assign v_RD_SIG11_3498_out0 = v_RD_SIG11_4356_out0;
assign v_Q_5096_out0 = v_OP2_SIG11_8_out0;
assign v_Q_5097_out0 = v_RD_SIG11_4356_out0;
assign v__5307_out0 = { v__2311_out0,v_G12_2294_out0 };
assign v_IN_6557_out0 = v_MUX2_1585_out0;
assign v__1407_out0 = v_IN_6557_out0[0:0];
assign v__1407_out1 = v_IN_6557_out0[15:15];
assign v__3753_out0 = { v_Q_5096_out0,v_C1_5084_out0 };
assign v__3754_out0 = { v_Q_5097_out0,v_C1_5085_out0 };
assign v__5079_out0 = { v__1584_out0,v_G6_6719_out0 };
assign v__5317_out0 = v_IN_6557_out0[15:15];
assign v_ADDER_IN_5411_out0 = v__5307_out0;
assign {v_A4_6704_out1,v_A4_6704_out0 } = v__5061_out0 + v_MUX8_2238_out0 + v_G4_6750_out0;
assign v__63_out0 = { v__5079_out0,v_G7_1357_out0 };
assign v__165_out0 = { v__1407_out1,v__5317_out0 };
assign v_UNUSED1_1472_out0 = v_A4_6704_out1;
assign v_NOTUSED_2183_out0 = v__1407_out0;
assign v_EXP_SUM_2864_out0 = v_A4_6704_out0;
assign v_OUT_3787_out0 = v__3753_out0;
assign v_OUT_3788_out0 = v__3754_out0;
assign v_SEL2_5089_out0 = v_A4_6704_out0[5:5];
assign v_RD_MULTI_25_out0 = v_OUT_3788_out0;
assign v_RM_MULTI_105_out0 = v_OUT_3787_out0;
assign {v_A6_1931_out1,v_A6_1931_out0 } = v_EXP_SUM_2864_out0 + v_MUX10_5120_out0 + v_0_5269_out0;
assign v_XOR4_3417_out0 = v_EXP_SUM_2864_out0 ^ v_NEG1_3398_out0;
assign v_OUT_5529_out0 = v__165_out0;
assign v_NEGATIVE_5541_out0 = v_SEL2_5089_out0;
assign v__6794_out0 = { v__63_out0,v_G8_596_out0 };
assign v_MUX4_137_out0 = v_NEGATIVE_5541_out0 ? v_OP2_EXP_5114_out0 : v_RD_EXP_1268_out0;
assign v__228_out0 = { v__6794_out0,v_G9_6552_out0 };
assign v_RM_MULTI_313_out0 = v_RM_MULTI_105_out0;
assign v_UNUSED2_1069_out0 = v_A6_1931_out1;
assign v_SHIFT_RD_1240_out0 = v_NEGATIVE_5541_out0;
assign {v_A5_1286_out1,v_A5_1286_out0 } = v_XOR4_3417_out0 + v_C11_6781_out0 + v_C10_888_out0;
assign v_RD_FLOATING_1379_out0 = v_RD_MULTI_25_out0;
assign v_SEL4_2837_out0 = v_A6_1931_out0[4:0];
assign v_MUX3_3474_out0 = v_ASR_4308_out0 ? v_OUT_5529_out0 : v_MUX2_1585_out0;
assign v_MUX11_46_out0 = v_G5_3486_out0 ? v_SEL4_2837_out0 : v_MUX4_137_out0;
assign v_UNUSED_168_out0 = v_A5_1286_out1;
assign v__207_out0 = { v__228_out0,v_G10_6518_out0 };
assign v_MUX7_572_out0 = v_FLOATING_INS_6796_out0 ? v_RD_FLOATING_1379_out0 : v_RD_245_out0;
assign v_MUX8_932_out0 = v_FLOATING_INS_6796_out0 ? v_RM_MULTI_313_out0 : v_RM_6773_out0;
assign v__1456_out0 = v_MUX3_3474_out0[0:0];
assign v__1456_out1 = v_MUX3_3474_out0[15:15];
assign v_G1_5295_out0 = ! v_SHIFT_RD_1240_out0;
assign v_MUX9_6643_out0 = v_NEGATIVE_5541_out0 ? v_A5_1286_out0 : v_EXP_SUM_2864_out0;
assign v_SEL3_190_out0 = v_MUX9_6643_out0[4:0];
assign v_RD_297_out0 = v_MUX7_572_out0;
assign v__1385_out0 = { v__207_out0,v_G11_6573_out0 };
assign v_RM_1591_out0 = v_MUX8_932_out0;
assign v__3492_out0 = { v__1456_out1,v__1456_out0 };
assign v_SHIFT_WHICH_OP_5274_out0 = v_G1_5295_out0;
assign v_EXP_ANS_5342_out0 = v_MUX11_46_out0;
assign v__212_out0 = v_RD_297_out0[2:2];
assign v__1314_out0 = v_RD_297_out0[1:1];
assign v_RM_1420_out0 = v_RM_1591_out0;
assign v__1550_out0 = v_RD_297_out0[3:3];
assign v_SHIFT_WHICH_OP_2181_out0 = v_SHIFT_WHICH_OP_5274_out0;
assign v_SHIFT_AMOUNT_2302_out0 = v_SEL3_190_out0;
assign v_RD_2362_out0 = v_RD_297_out0;
assign v_MUX4_3448_out0 = v_ROR_1599_out0 ? v__3492_out0 : v_MUX3_3474_out0;
assign v__3487_out0 = v_RD_297_out0[0:0];
assign v_A_5066_out0 = v_RM_1591_out0;
assign v_SHIFT_WHICH_OP_5153_out0 = v_SHIFT_WHICH_OP_5274_out0;
assign v_EXP_PRE_ANS_5299_out0 = v_EXP_ANS_5342_out0;
assign v_RM_5446_out0 = v_RM_1591_out0;
assign v_RM_5447_out0 = v_RM_1591_out0;
assign v_RM_5449_out0 = v_RM_1591_out0;
assign v__5483_out0 = { v__1385_out0,v_G12_1627_out0 };
assign v__0_out0 = v_A_5066_out0[4:4];
assign v__21_out0 = v_RD_2362_out0[7:7];
assign v_SHIFT_AMOUNT_113_out0 = v_SHIFT_AMOUNT_2302_out0;
assign v__247_out0 = v_RM_5446_out0[5:5];
assign v__248_out0 = v_RM_5447_out0[5:5];
assign v__250_out0 = v_RM_5449_out0[5:5];
assign v__278_out0 = v_RM_5446_out0[1:1];
assign v__279_out0 = v_RM_5447_out0[1:1];
assign v__281_out0 = v_RM_5449_out0[1:1];
assign v__577_out0 = v_RD_2362_out0[13:13];
assign v__584_out0 = v_RD_2362_out0[4:4];
assign v__831_out0 = v_A_5066_out0[5:5];
assign v__853_out0 = v_A_5066_out0[11:11];
assign v__926_out0 = v_A_5066_out0[0:0];
assign v__966_out0 = v_RM_5446_out0[15:15];
assign v__967_out0 = v_RM_5447_out0[15:15];
assign v__969_out0 = v_RM_5449_out0[15:15];
assign v__1008_out0 = v_RM_5446_out0[10:10];
assign v__1009_out0 = v_RM_5447_out0[10:10];
assign v__1011_out0 = v_RM_5449_out0[10:10];
assign v__1048_out0 = v_A_5066_out0[2:2];
assign v__1110_out0 = v_RM_5446_out0[12:12];
assign v__1111_out0 = v_RM_5447_out0[12:12];
assign v__1113_out0 = v_RM_5449_out0[12:12];
assign v_MUX1_1171_out0 = v_SHIFT_WHICH_OP_5153_out0 ? v__1352_out0 : v__3790_out0;
assign v__1203_out0 = v_RD_2362_out0[8:8];
assign v__1332_out0 = v_RM_5446_out0[2:2];
assign v__1333_out0 = v_RM_5447_out0[2:2];
assign v__1335_out0 = v_RM_5449_out0[2:2];
assign v__1347_out0 = v_A_5066_out0[15:15];
assign v__1401_out0 = v_A_5066_out0[12:12];
assign v__1403_out0 = v_A_5066_out0[3:3];
assign v_EXP_1416_out0 = v_EXP_PRE_ANS_5299_out0;
assign v__1451_out0 = v_RD_2362_out0[15:15];
assign v__1458_out0 = v_RM_5446_out0[8:8];
assign v__1459_out0 = v_RM_5447_out0[8:8];
assign v__1461_out0 = v_RM_5449_out0[8:8];
assign v__1558_out0 = { v__5483_out0,v_G13_2298_out0 };
assign v__1560_out0 = v_RD_2362_out0[10:10];
assign v__1580_out0 = v_A_5066_out0[8:8];
assign v_RDN_1628_out0 = v__3487_out0;
assign v__1854_out0 = v_RD_2362_out0[12:12];
assign v__1907_out0 = v_RM_5446_out0[11:11];
assign v__1908_out0 = v_RM_5447_out0[11:11];
assign v__1910_out0 = v_RM_5449_out0[11:11];
assign v__1934_out0 = v_RM_5446_out0[9:9];
assign v__1935_out0 = v_RM_5447_out0[9:9];
assign v__1937_out0 = v_RM_5449_out0[9:9];
assign v_RDN_2197_out0 = v__1314_out0;
assign v_RDN_2198_out0 = v__212_out0;
assign v_RDN_2200_out0 = v__1550_out0;
assign v__2244_out0 = v_A_5066_out0[10:10];
assign v__2300_out0 = v_A_5066_out0[13:13];
assign v__3356_out0 = v_RM_5446_out0[14:14];
assign v__3357_out0 = v_RM_5447_out0[14:14];
assign v__3359_out0 = v_RM_5449_out0[14:14];
assign v_MUX5_3445_out0 = v_EN_1136_out0 ? v_MUX4_3448_out0 : v_IN_6792_out0;
assign v__4353_out0 = v_A_5066_out0[14:14];
assign v__5128_out0 = v_RM_5446_out0[7:7];
assign v__5129_out0 = v_RM_5447_out0[7:7];
assign v__5131_out0 = v_RM_5449_out0[7:7];
assign v__5157_out0 = v_RD_2362_out0[9:9];
assign v__5160_out0 = v_RD_2362_out0[6:6];
assign v__5275_out0 = v_RD_2362_out0[14:14];
assign v__5350_out0 = v_RM_5446_out0[4:4];
assign v__5351_out0 = v_RM_5447_out0[4:4];
assign v__5353_out0 = v_RM_5449_out0[4:4];
assign v__5415_out0 = v_RM_5446_out0[0:0];
assign v__5416_out0 = v_RM_5447_out0[0:0];
assign v__5418_out0 = v_RM_5449_out0[0:0];
assign v_RM_5445_out0 = v_RM_1420_out0;
assign v_RM_5448_out0 = v_RM_1420_out0;
assign v_RM_5450_out0 = v_RM_1420_out0;
assign v_RM_5451_out0 = v_RM_1420_out0;
assign v_RM_5452_out0 = v_RM_1420_out0;
assign v_RM_5453_out0 = v_RM_1420_out0;
assign v_RM_5454_out0 = v_RM_1420_out0;
assign v_RM_5455_out0 = v_RM_1420_out0;
assign v_RM_5456_out0 = v_RM_1420_out0;
assign v_RM_5457_out0 = v_RM_1420_out0;
assign v_RM_5458_out0 = v_RM_1420_out0;
assign v_RM_5459_out0 = v_RM_1420_out0;
assign v__5464_out0 = v_RM_5446_out0[3:3];
assign v__5465_out0 = v_RM_5447_out0[3:3];
assign v__5467_out0 = v_RM_5449_out0[3:3];
assign v__5487_out0 = v_A_5066_out0[6:6];
assign v__6593_out0 = v_A_5066_out0[7:7];
assign v__6601_out0 = v_RM_5446_out0[6:6];
assign v__6602_out0 = v_RM_5447_out0[6:6];
assign v__6604_out0 = v_RM_5449_out0[6:6];
assign v__6618_out0 = v_RD_2362_out0[5:5];
assign v__6659_out0 = v_A_5066_out0[1:1];
assign v__6703_out0 = v_RD_2362_out0[11:11];
assign v__6714_out0 = v_A_5066_out0[9:9];
assign v__6757_out0 = v_RM_5446_out0[13:13];
assign v__6758_out0 = v_RM_5447_out0[13:13];
assign v__6760_out0 = v_RM_5449_out0[13:13];
assign v__90_out0 = { v__1558_out0,v_G14_2216_out0 };
assign v_G3_121_out0 = v_RDN_2197_out0 && v__1332_out0;
assign v_G3_122_out0 = v_RDN_2198_out0 && v__1333_out0;
assign v_G3_124_out0 = v_RDN_2200_out0 && v__1335_out0;
assign v_G4_170_out0 = v_RDN_2197_out0 && v__5464_out0;
assign v_G4_171_out0 = v_RDN_2198_out0 && v__5465_out0;
assign v_G4_173_out0 = v_RDN_2200_out0 && v__5467_out0;
assign v__246_out0 = v_RM_5445_out0[5:5];
assign v__249_out0 = v_RM_5448_out0[5:5];
assign v__251_out0 = v_RM_5450_out0[5:5];
assign v__252_out0 = v_RM_5451_out0[5:5];
assign v__253_out0 = v_RM_5452_out0[5:5];
assign v__254_out0 = v_RM_5453_out0[5:5];
assign v__255_out0 = v_RM_5454_out0[5:5];
assign v__256_out0 = v_RM_5455_out0[5:5];
assign v__257_out0 = v_RM_5456_out0[5:5];
assign v__258_out0 = v_RM_5457_out0[5:5];
assign v__259_out0 = v_RM_5458_out0[5:5];
assign v__260_out0 = v_RM_5459_out0[5:5];
assign v_G8_269_out0 = v__6593_out0 && v_RDN_1628_out0;
assign v__277_out0 = v_RM_5445_out0[1:1];
assign v__280_out0 = v_RM_5448_out0[1:1];
assign v__282_out0 = v_RM_5450_out0[1:1];
assign v__283_out0 = v_RM_5451_out0[1:1];
assign v__284_out0 = v_RM_5452_out0[1:1];
assign v__285_out0 = v_RM_5453_out0[1:1];
assign v__286_out0 = v_RM_5454_out0[1:1];
assign v__287_out0 = v_RM_5455_out0[1:1];
assign v__288_out0 = v_RM_5456_out0[1:1];
assign v__289_out0 = v_RM_5457_out0[1:1];
assign v__290_out0 = v_RM_5458_out0[1:1];
assign v__291_out0 = v_RM_5459_out0[1:1];
assign v_G14_298_out0 = v__2300_out0 && v_RDN_1628_out0;
assign v_G13_310_out0 = v__1401_out0 && v_RDN_1628_out0;
assign v_OUT_557_out0 = v_MUX5_3445_out0;
assign v_G2_884_out0 = v__6659_out0 && v_RDN_1628_out0;
assign v_G1_919_out0 = v__926_out0 && v_RDN_1628_out0;
assign v_G1_934_out0 = v_RDN_2197_out0 && v__278_out0;
assign v_G1_935_out0 = v_RDN_2198_out0 && v__279_out0;
assign v_G1_937_out0 = v_RDN_2200_out0 && v__281_out0;
assign v__965_out0 = v_RM_5445_out0[15:15];
assign v__968_out0 = v_RM_5448_out0[15:15];
assign v__970_out0 = v_RM_5450_out0[15:15];
assign v__971_out0 = v_RM_5451_out0[15:15];
assign v__972_out0 = v_RM_5452_out0[15:15];
assign v__973_out0 = v_RM_5453_out0[15:15];
assign v__974_out0 = v_RM_5454_out0[15:15];
assign v__975_out0 = v_RM_5455_out0[15:15];
assign v__976_out0 = v_RM_5456_out0[15:15];
assign v__977_out0 = v_RM_5457_out0[15:15];
assign v__978_out0 = v_RM_5458_out0[15:15];
assign v__979_out0 = v_RM_5459_out0[15:15];
assign v__1007_out0 = v_RM_5445_out0[10:10];
assign v__1010_out0 = v_RM_5448_out0[10:10];
assign v__1012_out0 = v_RM_5450_out0[10:10];
assign v__1013_out0 = v_RM_5451_out0[10:10];
assign v__1014_out0 = v_RM_5452_out0[10:10];
assign v__1015_out0 = v_RM_5453_out0[10:10];
assign v__1016_out0 = v_RM_5454_out0[10:10];
assign v__1017_out0 = v_RM_5455_out0[10:10];
assign v__1018_out0 = v_RM_5456_out0[10:10];
assign v__1019_out0 = v_RM_5457_out0[10:10];
assign v__1020_out0 = v_RM_5458_out0[10:10];
assign v__1021_out0 = v_RM_5459_out0[10:10];
assign v_G6_1031_out0 = v_RDN_2197_out0 && v__6601_out0;
assign v_G6_1032_out0 = v_RDN_2198_out0 && v__6602_out0;
assign v_G6_1034_out0 = v_RDN_2200_out0 && v__6604_out0;
assign v__1109_out0 = v_RM_5445_out0[12:12];
assign v__1112_out0 = v_RM_5448_out0[12:12];
assign v__1114_out0 = v_RM_5450_out0[12:12];
assign v__1115_out0 = v_RM_5451_out0[12:12];
assign v__1116_out0 = v_RM_5452_out0[12:12];
assign v__1117_out0 = v_RM_5453_out0[12:12];
assign v__1118_out0 = v_RM_5454_out0[12:12];
assign v__1119_out0 = v_RM_5455_out0[12:12];
assign v__1120_out0 = v_RM_5456_out0[12:12];
assign v__1121_out0 = v_RM_5457_out0[12:12];
assign v__1122_out0 = v_RM_5458_out0[12:12];
assign v__1123_out0 = v_RM_5459_out0[12:12];
assign v_EXP_1188_out0 = v_EXP_1416_out0;
assign v_G8_1206_out0 = v_RDN_2197_out0 && v__1458_out0;
assign v_G8_1207_out0 = v_RDN_2198_out0 && v__1459_out0;
assign v_G8_1209_out0 = v_RDN_2200_out0 && v__1461_out0;
assign v_G10_1287_out0 = v__6714_out0 && v_RDN_1628_out0;
assign v__1331_out0 = v_RM_5445_out0[2:2];
assign v__1334_out0 = v_RM_5448_out0[2:2];
assign v__1336_out0 = v_RM_5450_out0[2:2];
assign v__1337_out0 = v_RM_5451_out0[2:2];
assign v__1338_out0 = v_RM_5452_out0[2:2];
assign v__1339_out0 = v_RM_5453_out0[2:2];
assign v__1340_out0 = v_RM_5454_out0[2:2];
assign v__1341_out0 = v_RM_5455_out0[2:2];
assign v__1342_out0 = v_RM_5456_out0[2:2];
assign v__1343_out0 = v_RM_5457_out0[2:2];
assign v__1344_out0 = v_RM_5458_out0[2:2];
assign v__1345_out0 = v_RM_5459_out0[2:2];
assign v_G4_1350_out0 = v__1403_out0 && v_RDN_1628_out0;
assign v_G5_1358_out0 = v__0_out0 && v_RDN_1628_out0;
assign v_G9_1410_out0 = v__1580_out0 && v_RDN_1628_out0;
assign v_G11_1433_out0 = v__2244_out0 && v_RDN_1628_out0;
assign v__1457_out0 = v_RM_5445_out0[8:8];
assign v__1460_out0 = v_RM_5448_out0[8:8];
assign v__1462_out0 = v_RM_5450_out0[8:8];
assign v__1463_out0 = v_RM_5451_out0[8:8];
assign v__1464_out0 = v_RM_5452_out0[8:8];
assign v__1465_out0 = v_RM_5453_out0[8:8];
assign v__1466_out0 = v_RM_5454_out0[8:8];
assign v__1467_out0 = v_RM_5455_out0[8:8];
assign v__1468_out0 = v_RM_5456_out0[8:8];
assign v__1469_out0 = v_RM_5457_out0[8:8];
assign v__1470_out0 = v_RM_5458_out0[8:8];
assign v__1471_out0 = v_RM_5459_out0[8:8];
assign v__1906_out0 = v_RM_5445_out0[11:11];
assign v__1909_out0 = v_RM_5448_out0[11:11];
assign v__1911_out0 = v_RM_5450_out0[11:11];
assign v__1912_out0 = v_RM_5451_out0[11:11];
assign v__1913_out0 = v_RM_5452_out0[11:11];
assign v__1914_out0 = v_RM_5453_out0[11:11];
assign v__1915_out0 = v_RM_5454_out0[11:11];
assign v__1916_out0 = v_RM_5455_out0[11:11];
assign v__1917_out0 = v_RM_5456_out0[11:11];
assign v__1918_out0 = v_RM_5457_out0[11:11];
assign v__1919_out0 = v_RM_5458_out0[11:11];
assign v__1920_out0 = v_RM_5459_out0[11:11];
assign v_B_1924_out0 = v_SHIFT_AMOUNT_113_out0;
assign v__1933_out0 = v_RM_5445_out0[9:9];
assign v__1936_out0 = v_RM_5448_out0[9:9];
assign v__1938_out0 = v_RM_5450_out0[9:9];
assign v__1939_out0 = v_RM_5451_out0[9:9];
assign v__1940_out0 = v_RM_5452_out0[9:9];
assign v__1941_out0 = v_RM_5453_out0[9:9];
assign v__1942_out0 = v_RM_5454_out0[9:9];
assign v__1943_out0 = v_RM_5455_out0[9:9];
assign v__1944_out0 = v_RM_5456_out0[9:9];
assign v__1945_out0 = v_RM_5457_out0[9:9];
assign v__1946_out0 = v_RM_5458_out0[9:9];
assign v__1947_out0 = v_RM_5459_out0[9:9];
assign v_RDN_2196_out0 = v__584_out0;
assign v_RDN_2199_out0 = v__6703_out0;
assign v_RDN_2201_out0 = v__1560_out0;
assign v_RDN_2202_out0 = v__1451_out0;
assign v_RDN_2203_out0 = v__5275_out0;
assign v_RDN_2204_out0 = v__1854_out0;
assign v_RDN_2205_out0 = v__1203_out0;
assign v_RDN_2206_out0 = v__6618_out0;
assign v_RDN_2207_out0 = v__21_out0;
assign v_RDN_2208_out0 = v__577_out0;
assign v_RDN_2209_out0 = v__5160_out0;
assign v_RDN_2210_out0 = v__5157_out0;
assign v_G2_2258_out0 = v_RDN_2197_out0 && v__5350_out0;
assign v_G2_2259_out0 = v_RDN_2198_out0 && v__5351_out0;
assign v_G2_2261_out0 = v_RDN_2200_out0 && v__5353_out0;
assign v_G15_2274_out0 = v__4353_out0 && v_RDN_1628_out0;
assign v__3355_out0 = v_RM_5445_out0[14:14];
assign v__3358_out0 = v_RM_5448_out0[14:14];
assign v__3360_out0 = v_RM_5450_out0[14:14];
assign v__3361_out0 = v_RM_5451_out0[14:14];
assign v__3362_out0 = v_RM_5452_out0[14:14];
assign v__3363_out0 = v_RM_5453_out0[14:14];
assign v__3364_out0 = v_RM_5454_out0[14:14];
assign v__3365_out0 = v_RM_5455_out0[14:14];
assign v__3366_out0 = v_RM_5456_out0[14:14];
assign v__3367_out0 = v_RM_5457_out0[14:14];
assign v__3368_out0 = v_RM_5458_out0[14:14];
assign v__3369_out0 = v_RM_5459_out0[14:14];
assign v_EQ1_3415_out0 = v_EXP_1416_out0 == 5'h0;
assign v_G3_3479_out0 = v__1048_out0 && v_RDN_1628_out0;
assign v_G7_4260_out0 = v__5487_out0 && v_RDN_1628_out0;
assign v_G6_4346_out0 = v__831_out0 && v_RDN_1628_out0;
assign v__5127_out0 = v_RM_5445_out0[7:7];
assign v__5130_out0 = v_RM_5448_out0[7:7];
assign v__5132_out0 = v_RM_5450_out0[7:7];
assign v__5133_out0 = v_RM_5451_out0[7:7];
assign v__5134_out0 = v_RM_5452_out0[7:7];
assign v__5135_out0 = v_RM_5453_out0[7:7];
assign v__5136_out0 = v_RM_5454_out0[7:7];
assign v__5137_out0 = v_RM_5455_out0[7:7];
assign v__5138_out0 = v_RM_5456_out0[7:7];
assign v__5139_out0 = v_RM_5457_out0[7:7];
assign v__5140_out0 = v_RM_5458_out0[7:7];
assign v__5141_out0 = v_RM_5459_out0[7:7];
assign v_G9_5204_out0 = v_RDN_2197_out0 && v__1934_out0;
assign v_G9_5205_out0 = v_RDN_2198_out0 && v__1935_out0;
assign v_G9_5207_out0 = v_RDN_2200_out0 && v__1937_out0;
assign v_G5_5229_out0 = v_RDN_2197_out0 && v__247_out0;
assign v_G5_5230_out0 = v_RDN_2198_out0 && v__248_out0;
assign v_G5_5232_out0 = v_RDN_2200_out0 && v__250_out0;
assign v_G12_5261_out0 = v__853_out0 && v_RDN_1628_out0;
assign v_SIG_TO_SHIFT_5273_out0 = v_MUX1_1171_out0;
assign v__5349_out0 = v_RM_5445_out0[4:4];
assign v__5352_out0 = v_RM_5448_out0[4:4];
assign v__5354_out0 = v_RM_5450_out0[4:4];
assign v__5355_out0 = v_RM_5451_out0[4:4];
assign v__5356_out0 = v_RM_5452_out0[4:4];
assign v__5357_out0 = v_RM_5453_out0[4:4];
assign v__5358_out0 = v_RM_5454_out0[4:4];
assign v__5359_out0 = v_RM_5455_out0[4:4];
assign v__5360_out0 = v_RM_5456_out0[4:4];
assign v__5361_out0 = v_RM_5457_out0[4:4];
assign v__5362_out0 = v_RM_5458_out0[4:4];
assign v__5363_out0 = v_RM_5459_out0[4:4];
assign v_G16_5365_out0 = v__1347_out0 && v_RDN_1628_out0;
assign v__5414_out0 = v_RM_5445_out0[0:0];
assign v__5417_out0 = v_RM_5448_out0[0:0];
assign v__5419_out0 = v_RM_5450_out0[0:0];
assign v__5420_out0 = v_RM_5451_out0[0:0];
assign v__5421_out0 = v_RM_5452_out0[0:0];
assign v__5422_out0 = v_RM_5453_out0[0:0];
assign v__5423_out0 = v_RM_5454_out0[0:0];
assign v__5424_out0 = v_RM_5455_out0[0:0];
assign v__5425_out0 = v_RM_5456_out0[0:0];
assign v__5426_out0 = v_RM_5457_out0[0:0];
assign v__5427_out0 = v_RM_5458_out0[0:0];
assign v__5428_out0 = v_RM_5459_out0[0:0];
assign v__5463_out0 = v_RM_5445_out0[3:3];
assign v__5466_out0 = v_RM_5448_out0[3:3];
assign v__5468_out0 = v_RM_5450_out0[3:3];
assign v__5469_out0 = v_RM_5451_out0[3:3];
assign v__5470_out0 = v_RM_5452_out0[3:3];
assign v__5471_out0 = v_RM_5453_out0[3:3];
assign v__5472_out0 = v_RM_5454_out0[3:3];
assign v__5473_out0 = v_RM_5455_out0[3:3];
assign v__5474_out0 = v_RM_5456_out0[3:3];
assign v__5475_out0 = v_RM_5457_out0[3:3];
assign v__5476_out0 = v_RM_5458_out0[3:3];
assign v__5477_out0 = v_RM_5459_out0[3:3];
assign v_EQ2_5540_out0 = v_EXP_1416_out0 == 5'h1;
assign v_G7_5544_out0 = v_RDN_2197_out0 && v__5128_out0;
assign v_G7_5545_out0 = v_RDN_2198_out0 && v__5129_out0;
assign v_G7_5547_out0 = v_RDN_2200_out0 && v__5131_out0;
assign v_G16_6502_out0 = v_RDN_2197_out0 && v__5415_out0;
assign v_G16_6503_out0 = v_RDN_2198_out0 && v__5416_out0;
assign v_G16_6505_out0 = v_RDN_2200_out0 && v__5418_out0;
assign v__6600_out0 = v_RM_5445_out0[6:6];
assign v__6603_out0 = v_RM_5448_out0[6:6];
assign v__6605_out0 = v_RM_5450_out0[6:6];
assign v__6606_out0 = v_RM_5451_out0[6:6];
assign v__6607_out0 = v_RM_5452_out0[6:6];
assign v__6608_out0 = v_RM_5453_out0[6:6];
assign v__6609_out0 = v_RM_5454_out0[6:6];
assign v__6610_out0 = v_RM_5455_out0[6:6];
assign v__6611_out0 = v_RM_5456_out0[6:6];
assign v__6612_out0 = v_RM_5457_out0[6:6];
assign v__6613_out0 = v_RM_5458_out0[6:6];
assign v__6614_out0 = v_RM_5459_out0[6:6];
assign v_RD_6687_out0 = v_RDN_2197_out0;
assign v_RD_6688_out0 = v_RDN_2198_out0;
assign v_RD_6690_out0 = v_RDN_2200_out0;
assign v__6756_out0 = v_RM_5445_out0[13:13];
assign v__6759_out0 = v_RM_5448_out0[13:13];
assign v__6761_out0 = v_RM_5450_out0[13:13];
assign v__6762_out0 = v_RM_5451_out0[13:13];
assign v__6763_out0 = v_RM_5452_out0[13:13];
assign v__6764_out0 = v_RM_5453_out0[13:13];
assign v__6765_out0 = v_RM_5454_out0[13:13];
assign v__6766_out0 = v_RM_5455_out0[13:13];
assign v__6767_out0 = v_RM_5456_out0[13:13];
assign v__6768_out0 = v_RM_5457_out0[13:13];
assign v__6769_out0 = v_RM_5458_out0[13:13];
assign v__6770_out0 = v_RM_5459_out0[13:13];
assign v_G15_69_out0 = v_RD_6687_out0 && v__966_out0;
assign v_G15_70_out0 = v_RD_6688_out0 && v__967_out0;
assign v_G15_72_out0 = v_RD_6690_out0 && v__969_out0;
assign v_G3_120_out0 = v_RDN_2196_out0 && v__1331_out0;
assign v_G3_123_out0 = v_RDN_2199_out0 && v__1334_out0;
assign v_G3_125_out0 = v_RDN_2201_out0 && v__1336_out0;
assign v_G3_126_out0 = v_RDN_2202_out0 && v__1337_out0;
assign v_G3_127_out0 = v_RDN_2203_out0 && v__1338_out0;
assign v_G3_128_out0 = v_RDN_2204_out0 && v__1339_out0;
assign v_G3_129_out0 = v_RDN_2205_out0 && v__1340_out0;
assign v_G3_130_out0 = v_RDN_2206_out0 && v__1341_out0;
assign v_G3_131_out0 = v_RDN_2207_out0 && v__1342_out0;
assign v_G3_132_out0 = v_RDN_2208_out0 && v__1343_out0;
assign v_G3_133_out0 = v_RDN_2209_out0 && v__1344_out0;
assign v_G3_134_out0 = v_RDN_2210_out0 && v__1345_out0;
assign v_G4_169_out0 = v_RDN_2196_out0 && v__5463_out0;
assign v_G4_172_out0 = v_RDN_2199_out0 && v__5466_out0;
assign v_G4_174_out0 = v_RDN_2201_out0 && v__5468_out0;
assign v_G4_175_out0 = v_RDN_2202_out0 && v__5469_out0;
assign v_G4_176_out0 = v_RDN_2203_out0 && v__5470_out0;
assign v_G4_177_out0 = v_RDN_2204_out0 && v__5471_out0;
assign v_G4_178_out0 = v_RDN_2205_out0 && v__5472_out0;
assign v_G4_179_out0 = v_RDN_2206_out0 && v__5473_out0;
assign v_G4_180_out0 = v_RDN_2207_out0 && v__5474_out0;
assign v_G4_181_out0 = v_RDN_2208_out0 && v__5475_out0;
assign v_G4_182_out0 = v_RDN_2209_out0 && v__5476_out0;
assign v_G4_183_out0 = v_RDN_2210_out0 && v__5477_out0;
assign v__188_out0 = { v_G5_1358_out0,v_G6_4346_out0 };
assign v__193_out0 = { v_G9_1410_out0,v_G10_1287_out0 };
assign v_G11_316_out0 = v_RD_6687_out0 && v__1907_out0;
assign v_G11_317_out0 = v_RD_6688_out0 && v__1908_out0;
assign v_G11_319_out0 = v_RD_6690_out0 && v__1910_out0;
assign v_2_862_out0 = v_B_1924_out0[2:2];
assign v_G1_933_out0 = v_RDN_2196_out0 && v__277_out0;
assign v_G1_936_out0 = v_RDN_2199_out0 && v__280_out0;
assign v_G1_938_out0 = v_RDN_2201_out0 && v__282_out0;
assign v_G1_939_out0 = v_RDN_2202_out0 && v__283_out0;
assign v_G1_940_out0 = v_RDN_2203_out0 && v__284_out0;
assign v_G1_941_out0 = v_RDN_2204_out0 && v__285_out0;
assign v_G1_942_out0 = v_RDN_2205_out0 && v__286_out0;
assign v_G1_943_out0 = v_RDN_2206_out0 && v__287_out0;
assign v_G1_944_out0 = v_RDN_2207_out0 && v__288_out0;
assign v_G1_945_out0 = v_RDN_2208_out0 && v__289_out0;
assign v_G1_946_out0 = v_RDN_2209_out0 && v__290_out0;
assign v_G1_947_out0 = v_RDN_2210_out0 && v__291_out0;
assign v_G6_1030_out0 = v_RDN_2196_out0 && v__6600_out0;
assign v_G6_1033_out0 = v_RDN_2199_out0 && v__6603_out0;
assign v_G6_1035_out0 = v_RDN_2201_out0 && v__6605_out0;
assign v_G6_1036_out0 = v_RDN_2202_out0 && v__6606_out0;
assign v_G6_1037_out0 = v_RDN_2203_out0 && v__6607_out0;
assign v_G6_1038_out0 = v_RDN_2204_out0 && v__6608_out0;
assign v_G6_1039_out0 = v_RDN_2205_out0 && v__6609_out0;
assign v_G6_1040_out0 = v_RDN_2206_out0 && v__6610_out0;
assign v_G6_1041_out0 = v_RDN_2207_out0 && v__6611_out0;
assign v_G6_1042_out0 = v_RDN_2208_out0 && v__6612_out0;
assign v_G6_1043_out0 = v_RDN_2209_out0 && v__6613_out0;
assign v_G6_1044_out0 = v_RDN_2210_out0 && v__6614_out0;
assign v_G8_1205_out0 = v_RDN_2196_out0 && v__1457_out0;
assign v_G8_1208_out0 = v_RDN_2199_out0 && v__1460_out0;
assign v_G8_1210_out0 = v_RDN_2201_out0 && v__1462_out0;
assign v_G8_1211_out0 = v_RDN_2202_out0 && v__1463_out0;
assign v_G8_1212_out0 = v_RDN_2203_out0 && v__1464_out0;
assign v_G8_1213_out0 = v_RDN_2204_out0 && v__1465_out0;
assign v_G8_1214_out0 = v_RDN_2205_out0 && v__1466_out0;
assign v_G8_1215_out0 = v_RDN_2206_out0 && v__1467_out0;
assign v_G8_1216_out0 = v_RDN_2207_out0 && v__1468_out0;
assign v_G8_1217_out0 = v_RDN_2208_out0 && v__1469_out0;
assign v_G8_1218_out0 = v_RDN_2209_out0 && v__1470_out0;
assign v_G8_1219_out0 = v_RDN_2210_out0 && v__1471_out0;
assign v__1437_out0 = { v_G15_2274_out0,v_G16_5365_out0 };
assign v_0_1475_out0 = v_B_1924_out0[0:0];
assign v__1566_out0 = { v_G1_919_out0,v_G2_884_out0 };
assign v__1594_out0 = { v_G3_3479_out0,v_G4_1350_out0 };
assign v_1_1860_out0 = v_B_1924_out0[1:1];
assign v_G2_2257_out0 = v_RDN_2196_out0 && v__5349_out0;
assign v_G2_2260_out0 = v_RDN_2199_out0 && v__5352_out0;
assign v_G2_2262_out0 = v_RDN_2201_out0 && v__5354_out0;
assign v_G2_2263_out0 = v_RDN_2202_out0 && v__5355_out0;
assign v_G2_2264_out0 = v_RDN_2203_out0 && v__5356_out0;
assign v_G2_2265_out0 = v_RDN_2204_out0 && v__5357_out0;
assign v_G2_2266_out0 = v_RDN_2205_out0 && v__5358_out0;
assign v_G2_2267_out0 = v_RDN_2206_out0 && v__5359_out0;
assign v_G2_2268_out0 = v_RDN_2207_out0 && v__5360_out0;
assign v_G2_2269_out0 = v_RDN_2208_out0 && v__5361_out0;
assign v_G2_2270_out0 = v_RDN_2209_out0 && v__5362_out0;
assign v_G2_2271_out0 = v_RDN_2210_out0 && v__5363_out0;
assign v_SIG_TO_SHIFT_2861_out0 = v_SIG_TO_SHIFT_5273_out0;
assign v_RD_2913_out0 = v_G16_6502_out0;
assign v_RD_2945_out0 = v_G16_6503_out0;
assign v_RD_3007_out0 = v_G16_6505_out0;
assign v_G10_3425_out0 = v_RD_6687_out0 && v__1008_out0;
assign v_G10_3426_out0 = v_RD_6688_out0 && v__1009_out0;
assign v_G10_3428_out0 = v_RD_6690_out0 && v__1011_out0;
assign v__3501_out0 = { v_G13_310_out0,v_G14_298_out0 };
assign v_RD_3544_out0 = v_G5_5229_out0;
assign v_RD_3545_out0 = v_G2_2258_out0;
assign v_RD_3547_out0 = v_G9_5204_out0;
assign v_RD_3549_out0 = v_G1_934_out0;
assign v_RD_3550_out0 = v_G4_170_out0;
assign v_RD_3551_out0 = v_G6_1031_out0;
assign v_RD_3552_out0 = v_G7_5544_out0;
assign v_RD_3554_out0 = v_G8_1206_out0;
assign v_RD_3555_out0 = v_G3_121_out0;
assign v_RD_3559_out0 = v_G5_5230_out0;
assign v_RD_3560_out0 = v_G2_2259_out0;
assign v_RD_3562_out0 = v_G9_5205_out0;
assign v_RD_3564_out0 = v_G1_935_out0;
assign v_RD_3565_out0 = v_G4_171_out0;
assign v_RD_3566_out0 = v_G6_1032_out0;
assign v_RD_3567_out0 = v_G7_5545_out0;
assign v_RD_3569_out0 = v_G8_1207_out0;
assign v_RD_3570_out0 = v_G3_122_out0;
assign v_RD_3589_out0 = v_G5_5232_out0;
assign v_RD_3590_out0 = v_G2_2261_out0;
assign v_RD_3592_out0 = v_G9_5207_out0;
assign v_RD_3594_out0 = v_G1_937_out0;
assign v_RD_3595_out0 = v_G4_173_out0;
assign v_RD_3596_out0 = v_G6_1034_out0;
assign v_RD_3597_out0 = v_G7_5547_out0;
assign v_RD_3599_out0 = v_G8_1209_out0;
assign v_RD_3600_out0 = v_G3_124_out0;
assign v_SUBNORMAL_4335_out0 = v_EQ1_3415_out0;
assign v_IN_5124_out0 = v_OUT_557_out0;
assign v__5150_out0 = { v__90_out0,v_G15_887_out0 };
assign v_G9_5203_out0 = v_RDN_2196_out0 && v__1933_out0;
assign v_G9_5206_out0 = v_RDN_2199_out0 && v__1936_out0;
assign v_G9_5208_out0 = v_RDN_2201_out0 && v__1938_out0;
assign v_G9_5209_out0 = v_RDN_2202_out0 && v__1939_out0;
assign v_G9_5210_out0 = v_RDN_2203_out0 && v__1940_out0;
assign v_G9_5211_out0 = v_RDN_2204_out0 && v__1941_out0;
assign v_G9_5212_out0 = v_RDN_2205_out0 && v__1942_out0;
assign v_G9_5213_out0 = v_RDN_2206_out0 && v__1943_out0;
assign v_G9_5214_out0 = v_RDN_2207_out0 && v__1944_out0;
assign v_G9_5215_out0 = v_RDN_2208_out0 && v__1945_out0;
assign v_G9_5216_out0 = v_RDN_2209_out0 && v__1946_out0;
assign v_G9_5217_out0 = v_RDN_2210_out0 && v__1947_out0;
assign v_G5_5228_out0 = v_RDN_2196_out0 && v__246_out0;
assign v_G5_5231_out0 = v_RDN_2199_out0 && v__249_out0;
assign v_G5_5233_out0 = v_RDN_2201_out0 && v__251_out0;
assign v_G5_5234_out0 = v_RDN_2202_out0 && v__252_out0;
assign v_G5_5235_out0 = v_RDN_2203_out0 && v__253_out0;
assign v_G5_5236_out0 = v_RDN_2204_out0 && v__254_out0;
assign v_G5_5237_out0 = v_RDN_2205_out0 && v__255_out0;
assign v_G5_5238_out0 = v_RDN_2206_out0 && v__256_out0;
assign v_G5_5239_out0 = v_RDN_2207_out0 && v__257_out0;
assign v_G5_5240_out0 = v_RDN_2208_out0 && v__258_out0;
assign v_G5_5241_out0 = v_RDN_2209_out0 && v__259_out0;
assign v_G5_5242_out0 = v_RDN_2210_out0 && v__260_out0;
assign v_G7_5543_out0 = v_RDN_2196_out0 && v__5127_out0;
assign v_G7_5546_out0 = v_RDN_2199_out0 && v__5130_out0;
assign v_G7_5548_out0 = v_RDN_2201_out0 && v__5132_out0;
assign v_G7_5549_out0 = v_RDN_2202_out0 && v__5133_out0;
assign v_G7_5550_out0 = v_RDN_2203_out0 && v__5134_out0;
assign v_G7_5551_out0 = v_RDN_2204_out0 && v__5135_out0;
assign v_G7_5552_out0 = v_RDN_2205_out0 && v__5136_out0;
assign v_G7_5553_out0 = v_RDN_2206_out0 && v__5137_out0;
assign v_G7_5554_out0 = v_RDN_2207_out0 && v__5138_out0;
assign v_G7_5555_out0 = v_RDN_2208_out0 && v__5139_out0;
assign v_G7_5556_out0 = v_RDN_2209_out0 && v__5140_out0;
assign v_G7_5557_out0 = v_RDN_2210_out0 && v__5141_out0;
assign v_G16_6501_out0 = v_RDN_2196_out0 && v__5414_out0;
assign v_G16_6504_out0 = v_RDN_2199_out0 && v__5417_out0;
assign v_G16_6506_out0 = v_RDN_2201_out0 && v__5419_out0;
assign v_G16_6507_out0 = v_RDN_2202_out0 && v__5420_out0;
assign v_G16_6508_out0 = v_RDN_2203_out0 && v__5421_out0;
assign v_G16_6509_out0 = v_RDN_2204_out0 && v__5422_out0;
assign v_G16_6510_out0 = v_RDN_2205_out0 && v__5423_out0;
assign v_G16_6511_out0 = v_RDN_2206_out0 && v__5424_out0;
assign v_G16_6512_out0 = v_RDN_2207_out0 && v__5425_out0;
assign v_G16_6513_out0 = v_RDN_2208_out0 && v__5426_out0;
assign v_G16_6514_out0 = v_RDN_2209_out0 && v__5427_out0;
assign v_G16_6515_out0 = v_RDN_2210_out0 && v__5428_out0;
assign v_G12_6521_out0 = v_RD_6687_out0 && v__1110_out0;
assign v_G12_6522_out0 = v_RD_6688_out0 && v__1111_out0;
assign v_G12_6524_out0 = v_RD_6690_out0 && v__1113_out0;
assign v__6538_out0 = { v_G11_1433_out0,v_G12_5261_out0 };
assign v_G13_6578_out0 = v_RD_6687_out0 && v__6757_out0;
assign v_G13_6579_out0 = v_RD_6688_out0 && v__6758_out0;
assign v_G13_6581_out0 = v_RD_6690_out0 && v__6760_out0;
assign v_EXP1_6644_out0 = v_EQ2_5540_out0;
assign v_RD_6686_out0 = v_RDN_2196_out0;
assign v_RD_6689_out0 = v_RDN_2199_out0;
assign v_RD_6691_out0 = v_RDN_2201_out0;
assign v_RD_6692_out0 = v_RDN_2202_out0;
assign v_RD_6693_out0 = v_RDN_2203_out0;
assign v_RD_6694_out0 = v_RDN_2204_out0;
assign v_RD_6695_out0 = v_RDN_2205_out0;
assign v_RD_6696_out0 = v_RDN_2206_out0;
assign v_RD_6697_out0 = v_RDN_2207_out0;
assign v_RD_6698_out0 = v_RDN_2208_out0;
assign v_RD_6699_out0 = v_RDN_2209_out0;
assign v_RD_6700_out0 = v_RDN_2210_out0;
assign v_3_6711_out0 = v_B_1924_out0[3:3];
assign v_G14_6736_out0 = v_RD_6687_out0 && v__3356_out0;
assign v_G14_6737_out0 = v_RD_6688_out0 && v__3357_out0;
assign v_G14_6739_out0 = v_RD_6690_out0 && v__3359_out0;
assign v__6783_out0 = { v_G7_4260_out0,v_G8_269_out0 };
assign v__59_out0 = { v__188_out0,v__6783_out0 };
assign v_G15_68_out0 = v_RD_6686_out0 && v__965_out0;
assign v_G15_71_out0 = v_RD_6689_out0 && v__968_out0;
assign v_G15_73_out0 = v_RD_6691_out0 && v__970_out0;
assign v_G15_74_out0 = v_RD_6692_out0 && v__971_out0;
assign v_G15_75_out0 = v_RD_6693_out0 && v__972_out0;
assign v_G15_76_out0 = v_RD_6694_out0 && v__973_out0;
assign v_G15_77_out0 = v_RD_6695_out0 && v__974_out0;
assign v_G15_78_out0 = v_RD_6696_out0 && v__975_out0;
assign v_G15_79_out0 = v_RD_6697_out0 && v__976_out0;
assign v_G15_80_out0 = v_RD_6698_out0 && v__977_out0;
assign v_G15_81_out0 = v_RD_6699_out0 && v__978_out0;
assign v_G15_82_out0 = v_RD_6700_out0 && v__979_out0;
assign v__219_out0 = { v__3501_out0,v__1437_out0 };
assign v_G5_309_out0 = ! v_EXP1_6644_out0;
assign v_G11_315_out0 = v_RD_6686_out0 && v__1906_out0;
assign v_G11_318_out0 = v_RD_6689_out0 && v__1909_out0;
assign v_G11_320_out0 = v_RD_6691_out0 && v__1911_out0;
assign v_G11_321_out0 = v_RD_6692_out0 && v__1912_out0;
assign v_G11_322_out0 = v_RD_6693_out0 && v__1913_out0;
assign v_G11_323_out0 = v_RD_6694_out0 && v__1914_out0;
assign v_G11_324_out0 = v_RD_6695_out0 && v__1915_out0;
assign v_G11_325_out0 = v_RD_6696_out0 && v__1916_out0;
assign v_G11_326_out0 = v_RD_6697_out0 && v__1917_out0;
assign v_G11_327_out0 = v_RD_6698_out0 && v__1918_out0;
assign v_G11_328_out0 = v_RD_6699_out0 && v__1919_out0;
assign v_G11_329_out0 = v_RD_6700_out0 && v__1920_out0;
assign v__594_out0 = { v__5150_out0,v_G16_5431_out0 };
assign v__1143_out0 = { v__193_out0,v__6538_out0 };
assign v_RD_2884_out0 = v_G16_6501_out0;
assign v_RD_2907_out0 = v_RD_3544_out0;
assign v_RD_2909_out0 = v_RD_3545_out0;
assign v_RD_2914_out0 = v_G15_69_out0;
assign v_RD_2915_out0 = v_RD_3547_out0;
assign v_RD_2919_out0 = v_RD_3549_out0;
assign v_RD_2921_out0 = v_RD_3550_out0;
assign v_RD_2923_out0 = v_RD_3551_out0;
assign v_RD_2925_out0 = v_RD_3552_out0;
assign v_RD_2929_out0 = v_RD_3554_out0;
assign v_RD_2931_out0 = v_RD_3555_out0;
assign v_RD_2939_out0 = v_RD_3559_out0;
assign v_RD_2941_out0 = v_RD_3560_out0;
assign v_RD_2946_out0 = v_RD_3562_out0;
assign v_RD_2950_out0 = v_RD_3564_out0;
assign v_RD_2952_out0 = v_RD_3565_out0;
assign v_RD_2954_out0 = v_RD_3566_out0;
assign v_RD_2956_out0 = v_RD_3567_out0;
assign v_RD_2960_out0 = v_RD_3569_out0;
assign v_RD_2962_out0 = v_RD_3570_out0;
assign v_RD_2976_out0 = v_G16_6504_out0;
assign v_RD_3001_out0 = v_RD_3589_out0;
assign v_RD_3003_out0 = v_RD_3590_out0;
assign v_RD_3008_out0 = v_RD_3592_out0;
assign v_RD_3012_out0 = v_RD_3594_out0;
assign v_RD_3014_out0 = v_RD_3595_out0;
assign v_RD_3016_out0 = v_RD_3596_out0;
assign v_RD_3018_out0 = v_RD_3597_out0;
assign v_RD_3022_out0 = v_RD_3599_out0;
assign v_RD_3024_out0 = v_RD_3600_out0;
assign v_RD_3038_out0 = v_G16_6506_out0;
assign v_RD_3069_out0 = v_G16_6507_out0;
assign v_RD_3100_out0 = v_G16_6508_out0;
assign v_RD_3131_out0 = v_G16_6509_out0;
assign v_RD_3162_out0 = v_G16_6510_out0;
assign v_RD_3193_out0 = v_G16_6511_out0;
assign v_RD_3224_out0 = v_G16_6512_out0;
assign v_RD_3255_out0 = v_G16_6513_out0;
assign v_RD_3286_out0 = v_G16_6514_out0;
assign v_RD_3317_out0 = v_G16_6515_out0;
assign v_G10_3424_out0 = v_RD_6686_out0 && v__1007_out0;
assign v_G10_3427_out0 = v_RD_6689_out0 && v__1010_out0;
assign v_G10_3429_out0 = v_RD_6691_out0 && v__1012_out0;
assign v_G10_3430_out0 = v_RD_6692_out0 && v__1013_out0;
assign v_G10_3431_out0 = v_RD_6693_out0 && v__1014_out0;
assign v_G10_3432_out0 = v_RD_6694_out0 && v__1015_out0;
assign v_G10_3433_out0 = v_RD_6695_out0 && v__1016_out0;
assign v_G10_3434_out0 = v_RD_6696_out0 && v__1017_out0;
assign v_G10_3435_out0 = v_RD_6697_out0 && v__1018_out0;
assign v_G10_3436_out0 = v_RD_6698_out0 && v__1019_out0;
assign v_G10_3437_out0 = v_RD_6699_out0 && v__1020_out0;
assign v_G10_3438_out0 = v_RD_6700_out0 && v__1021_out0;
assign v_RD_3530_out0 = v_G5_5228_out0;
assign v_RD_3531_out0 = v_G2_2257_out0;
assign v_RD_3533_out0 = v_G9_5203_out0;
assign v_RD_3535_out0 = v_G1_933_out0;
assign v_RD_3536_out0 = v_G4_169_out0;
assign v_RD_3537_out0 = v_G6_1030_out0;
assign v_RD_3538_out0 = v_G7_5543_out0;
assign v_RD_3540_out0 = v_G8_1205_out0;
assign v_RD_3541_out0 = v_G3_120_out0;
assign v_RD_3542_out0 = v_G12_6521_out0;
assign v_RD_3543_out0 = v_G14_6736_out0;
assign v_RD_3546_out0 = v_G13_6578_out0;
assign v_RD_3548_out0 = v_G10_3425_out0;
assign v_RD_3553_out0 = v_G11_316_out0;
assign v_RD_3556_out0 = v_G12_6522_out0;
assign v_RD_3557_out0 = v_G14_6737_out0;
assign v_RD_3558_out0 = v_G15_70_out0;
assign v_RD_3561_out0 = v_G13_6579_out0;
assign v_RD_3563_out0 = v_G10_3426_out0;
assign v_RD_3568_out0 = v_G11_317_out0;
assign v_RD_3574_out0 = v_G5_5231_out0;
assign v_RD_3575_out0 = v_G2_2260_out0;
assign v_RD_3577_out0 = v_G9_5206_out0;
assign v_RD_3579_out0 = v_G1_936_out0;
assign v_RD_3580_out0 = v_G4_172_out0;
assign v_RD_3581_out0 = v_G6_1033_out0;
assign v_RD_3582_out0 = v_G7_5546_out0;
assign v_RD_3584_out0 = v_G8_1208_out0;
assign v_RD_3585_out0 = v_G3_123_out0;
assign v_RD_3586_out0 = v_G12_6524_out0;
assign v_RD_3587_out0 = v_G14_6739_out0;
assign v_RD_3588_out0 = v_G15_72_out0;
assign v_RD_3591_out0 = v_G13_6581_out0;
assign v_RD_3593_out0 = v_G10_3428_out0;
assign v_RD_3598_out0 = v_G11_319_out0;
assign v_RD_3604_out0 = v_G5_5233_out0;
assign v_RD_3605_out0 = v_G2_2262_out0;
assign v_RD_3607_out0 = v_G9_5208_out0;
assign v_RD_3609_out0 = v_G1_938_out0;
assign v_RD_3610_out0 = v_G4_174_out0;
assign v_RD_3611_out0 = v_G6_1035_out0;
assign v_RD_3612_out0 = v_G7_5548_out0;
assign v_RD_3614_out0 = v_G8_1210_out0;
assign v_RD_3615_out0 = v_G3_125_out0;
assign v_RD_3619_out0 = v_G5_5234_out0;
assign v_RD_3620_out0 = v_G2_2263_out0;
assign v_RD_3622_out0 = v_G9_5209_out0;
assign v_RD_3624_out0 = v_G1_939_out0;
assign v_RD_3625_out0 = v_G4_175_out0;
assign v_RD_3626_out0 = v_G6_1036_out0;
assign v_RD_3627_out0 = v_G7_5549_out0;
assign v_RD_3629_out0 = v_G8_1211_out0;
assign v_RD_3630_out0 = v_G3_126_out0;
assign v_RD_3634_out0 = v_G5_5235_out0;
assign v_RD_3635_out0 = v_G2_2264_out0;
assign v_RD_3637_out0 = v_G9_5210_out0;
assign v_RD_3639_out0 = v_G1_940_out0;
assign v_RD_3640_out0 = v_G4_176_out0;
assign v_RD_3641_out0 = v_G6_1037_out0;
assign v_RD_3642_out0 = v_G7_5550_out0;
assign v_RD_3644_out0 = v_G8_1212_out0;
assign v_RD_3645_out0 = v_G3_127_out0;
assign v_RD_3649_out0 = v_G5_5236_out0;
assign v_RD_3650_out0 = v_G2_2265_out0;
assign v_RD_3652_out0 = v_G9_5211_out0;
assign v_RD_3654_out0 = v_G1_941_out0;
assign v_RD_3655_out0 = v_G4_177_out0;
assign v_RD_3656_out0 = v_G6_1038_out0;
assign v_RD_3657_out0 = v_G7_5551_out0;
assign v_RD_3659_out0 = v_G8_1213_out0;
assign v_RD_3660_out0 = v_G3_128_out0;
assign v_RD_3664_out0 = v_G5_5237_out0;
assign v_RD_3665_out0 = v_G2_2266_out0;
assign v_RD_3667_out0 = v_G9_5212_out0;
assign v_RD_3669_out0 = v_G1_942_out0;
assign v_RD_3670_out0 = v_G4_178_out0;
assign v_RD_3671_out0 = v_G6_1039_out0;
assign v_RD_3672_out0 = v_G7_5552_out0;
assign v_RD_3674_out0 = v_G8_1214_out0;
assign v_RD_3675_out0 = v_G3_129_out0;
assign v_RD_3679_out0 = v_G5_5238_out0;
assign v_RD_3680_out0 = v_G2_2267_out0;
assign v_RD_3682_out0 = v_G9_5213_out0;
assign v_RD_3684_out0 = v_G1_943_out0;
assign v_RD_3685_out0 = v_G4_179_out0;
assign v_RD_3686_out0 = v_G6_1040_out0;
assign v_RD_3687_out0 = v_G7_5553_out0;
assign v_RD_3689_out0 = v_G8_1215_out0;
assign v_RD_3690_out0 = v_G3_130_out0;
assign v_RD_3694_out0 = v_G5_5239_out0;
assign v_RD_3695_out0 = v_G2_2268_out0;
assign v_RD_3697_out0 = v_G9_5214_out0;
assign v_RD_3699_out0 = v_G1_944_out0;
assign v_RD_3700_out0 = v_G4_180_out0;
assign v_RD_3701_out0 = v_G6_1041_out0;
assign v_RD_3702_out0 = v_G7_5554_out0;
assign v_RD_3704_out0 = v_G8_1216_out0;
assign v_RD_3705_out0 = v_G3_131_out0;
assign v_RD_3709_out0 = v_G5_5240_out0;
assign v_RD_3710_out0 = v_G2_2269_out0;
assign v_RD_3712_out0 = v_G9_5215_out0;
assign v_RD_3714_out0 = v_G1_945_out0;
assign v_RD_3715_out0 = v_G4_181_out0;
assign v_RD_3716_out0 = v_G6_1042_out0;
assign v_RD_3717_out0 = v_G7_5555_out0;
assign v_RD_3719_out0 = v_G8_1217_out0;
assign v_RD_3720_out0 = v_G3_132_out0;
assign v_RD_3724_out0 = v_G5_5241_out0;
assign v_RD_3725_out0 = v_G2_2270_out0;
assign v_RD_3727_out0 = v_G9_5216_out0;
assign v_RD_3729_out0 = v_G1_946_out0;
assign v_RD_3730_out0 = v_G4_182_out0;
assign v_RD_3731_out0 = v_G6_1043_out0;
assign v_RD_3732_out0 = v_G7_5556_out0;
assign v_RD_3734_out0 = v_G8_1218_out0;
assign v_RD_3735_out0 = v_G3_133_out0;
assign v_RD_3739_out0 = v_G5_5242_out0;
assign v_RD_3740_out0 = v_G2_2271_out0;
assign v_RD_3742_out0 = v_G9_5217_out0;
assign v_RD_3744_out0 = v_G1_947_out0;
assign v_RD_3745_out0 = v_G4_183_out0;
assign v_RD_3746_out0 = v_G6_1044_out0;
assign v_RD_3747_out0 = v_G7_5557_out0;
assign v_RD_3749_out0 = v_G8_1219_out0;
assign v_RD_3750_out0 = v_G3_134_out0;
assign v_IN_4348_out0 = v_IN_5124_out0;
assign v__5109_out0 = { v__1566_out0,v__1594_out0 };
assign v__5437_out0 = v_IN_5124_out0[13:0];
assign v__5437_out1 = v_IN_5124_out0[15:2];
assign v_G12_6520_out0 = v_RD_6686_out0 && v__1109_out0;
assign v_G12_6523_out0 = v_RD_6689_out0 && v__1112_out0;
assign v_G12_6525_out0 = v_RD_6691_out0 && v__1114_out0;
assign v_G12_6526_out0 = v_RD_6692_out0 && v__1115_out0;
assign v_G12_6527_out0 = v_RD_6693_out0 && v__1116_out0;
assign v_G12_6528_out0 = v_RD_6694_out0 && v__1117_out0;
assign v_G12_6529_out0 = v_RD_6695_out0 && v__1118_out0;
assign v_G12_6530_out0 = v_RD_6696_out0 && v__1119_out0;
assign v_G12_6531_out0 = v_RD_6697_out0 && v__1120_out0;
assign v_G12_6532_out0 = v_RD_6698_out0 && v__1121_out0;
assign v_G12_6533_out0 = v_RD_6699_out0 && v__1122_out0;
assign v_G12_6534_out0 = v_RD_6700_out0 && v__1123_out0;
assign v_G13_6577_out0 = v_RD_6686_out0 && v__6756_out0;
assign v_G13_6580_out0 = v_RD_6689_out0 && v__6759_out0;
assign v_G13_6582_out0 = v_RD_6691_out0 && v__6761_out0;
assign v_G13_6583_out0 = v_RD_6692_out0 && v__6762_out0;
assign v_G13_6584_out0 = v_RD_6693_out0 && v__6763_out0;
assign v_G13_6585_out0 = v_RD_6694_out0 && v__6764_out0;
assign v_G13_6586_out0 = v_RD_6695_out0 && v__6765_out0;
assign v_G13_6587_out0 = v_RD_6696_out0 && v__6766_out0;
assign v_G13_6588_out0 = v_RD_6697_out0 && v__6767_out0;
assign v_G13_6589_out0 = v_RD_6698_out0 && v__6768_out0;
assign v_G13_6590_out0 = v_RD_6699_out0 && v__6769_out0;
assign v_G13_6591_out0 = v_RD_6700_out0 && v__6770_out0;
assign v_IN_6733_out0 = v_SIG_TO_SHIFT_2861_out0;
assign v_G14_6735_out0 = v_RD_6686_out0 && v__3355_out0;
assign v_G14_6738_out0 = v_RD_6689_out0 && v__3358_out0;
assign v_G14_6740_out0 = v_RD_6691_out0 && v__3360_out0;
assign v_G14_6741_out0 = v_RD_6692_out0 && v__3361_out0;
assign v_G14_6742_out0 = v_RD_6693_out0 && v__3362_out0;
assign v_G14_6743_out0 = v_RD_6694_out0 && v__3363_out0;
assign v_G14_6744_out0 = v_RD_6695_out0 && v__3364_out0;
assign v_G14_6745_out0 = v_RD_6696_out0 && v__3365_out0;
assign v_G14_6746_out0 = v_RD_6697_out0 && v__3366_out0;
assign v_G14_6747_out0 = v_RD_6698_out0 && v__3367_out0;
assign v_G14_6748_out0 = v_RD_6699_out0 && v__3368_out0;
assign v_G14_6749_out0 = v_RD_6700_out0 && v__3369_out0;
assign v_IN1_1067_out0 = v_IN_6733_out0;
assign v_NOTUSED_1262_out0 = v__5437_out1;
assign v__1310_out0 = { v__5109_out0,v__59_out0 };
assign v__2176_out0 = { v__1143_out0,v__219_out0 };
assign v_RD_2878_out0 = v_RD_3530_out0;
assign v_RD_2880_out0 = v_RD_3531_out0;
assign v_RD_2885_out0 = v_RD_3533_out0;
assign v_RD_2889_out0 = v_RD_3535_out0;
assign v_RD_2891_out0 = v_RD_3536_out0;
assign v_RD_2893_out0 = v_RD_3537_out0;
assign v_RD_2895_out0 = v_RD_3538_out0;
assign v_RD_2899_out0 = v_RD_3540_out0;
assign v_RD_2901_out0 = v_RD_3541_out0;
assign v_RD_2903_out0 = v_RD_3542_out0;
assign v_RD_2905_out0 = v_RD_3543_out0;
assign v_RD_2911_out0 = v_RD_3546_out0;
assign v_RD_2917_out0 = v_RD_3548_out0;
assign v_RD_2927_out0 = v_RD_3553_out0;
assign v_RD_2933_out0 = v_RD_3556_out0;
assign v_RD_2935_out0 = v_RD_3557_out0;
assign v_RD_2937_out0 = v_RD_3558_out0;
assign v_RD_2943_out0 = v_RD_3561_out0;
assign v_RD_2948_out0 = v_RD_3563_out0;
assign v_RD_2958_out0 = v_RD_3568_out0;
assign v_RD_2970_out0 = v_RD_3574_out0;
assign v_RD_2972_out0 = v_RD_3575_out0;
assign v_RD_2977_out0 = v_RD_3577_out0;
assign v_RD_2981_out0 = v_RD_3579_out0;
assign v_RD_2983_out0 = v_RD_3580_out0;
assign v_RD_2985_out0 = v_RD_3581_out0;
assign v_RD_2987_out0 = v_RD_3582_out0;
assign v_RD_2991_out0 = v_RD_3584_out0;
assign v_RD_2993_out0 = v_RD_3585_out0;
assign v_RD_2995_out0 = v_RD_3586_out0;
assign v_RD_2997_out0 = v_RD_3587_out0;
assign v_RD_2999_out0 = v_RD_3588_out0;
assign v_RD_3005_out0 = v_RD_3591_out0;
assign v_RD_3010_out0 = v_RD_3593_out0;
assign v_RD_3020_out0 = v_RD_3598_out0;
assign v_RD_3032_out0 = v_RD_3604_out0;
assign v_RD_3034_out0 = v_RD_3605_out0;
assign v_RD_3039_out0 = v_RD_3607_out0;
assign v_RD_3043_out0 = v_RD_3609_out0;
assign v_RD_3045_out0 = v_RD_3610_out0;
assign v_RD_3047_out0 = v_RD_3611_out0;
assign v_RD_3049_out0 = v_RD_3612_out0;
assign v_RD_3053_out0 = v_RD_3614_out0;
assign v_RD_3055_out0 = v_RD_3615_out0;
assign v_RD_3063_out0 = v_RD_3619_out0;
assign v_RD_3065_out0 = v_RD_3620_out0;
assign v_RD_3070_out0 = v_RD_3622_out0;
assign v_RD_3074_out0 = v_RD_3624_out0;
assign v_RD_3076_out0 = v_RD_3625_out0;
assign v_RD_3078_out0 = v_RD_3626_out0;
assign v_RD_3080_out0 = v_RD_3627_out0;
assign v_RD_3084_out0 = v_RD_3629_out0;
assign v_RD_3086_out0 = v_RD_3630_out0;
assign v_RD_3094_out0 = v_RD_3634_out0;
assign v_RD_3096_out0 = v_RD_3635_out0;
assign v_RD_3101_out0 = v_RD_3637_out0;
assign v_RD_3105_out0 = v_RD_3639_out0;
assign v_RD_3107_out0 = v_RD_3640_out0;
assign v_RD_3109_out0 = v_RD_3641_out0;
assign v_RD_3111_out0 = v_RD_3642_out0;
assign v_RD_3115_out0 = v_RD_3644_out0;
assign v_RD_3117_out0 = v_RD_3645_out0;
assign v_RD_3125_out0 = v_RD_3649_out0;
assign v_RD_3127_out0 = v_RD_3650_out0;
assign v_RD_3132_out0 = v_RD_3652_out0;
assign v_RD_3136_out0 = v_RD_3654_out0;
assign v_RD_3138_out0 = v_RD_3655_out0;
assign v_RD_3140_out0 = v_RD_3656_out0;
assign v_RD_3142_out0 = v_RD_3657_out0;
assign v_RD_3146_out0 = v_RD_3659_out0;
assign v_RD_3148_out0 = v_RD_3660_out0;
assign v_RD_3156_out0 = v_RD_3664_out0;
assign v_RD_3158_out0 = v_RD_3665_out0;
assign v_RD_3163_out0 = v_RD_3667_out0;
assign v_RD_3167_out0 = v_RD_3669_out0;
assign v_RD_3169_out0 = v_RD_3670_out0;
assign v_RD_3171_out0 = v_RD_3671_out0;
assign v_RD_3173_out0 = v_RD_3672_out0;
assign v_RD_3177_out0 = v_RD_3674_out0;
assign v_RD_3179_out0 = v_RD_3675_out0;
assign v_RD_3187_out0 = v_RD_3679_out0;
assign v_RD_3189_out0 = v_RD_3680_out0;
assign v_RD_3194_out0 = v_RD_3682_out0;
assign v_RD_3198_out0 = v_RD_3684_out0;
assign v_RD_3200_out0 = v_RD_3685_out0;
assign v_RD_3202_out0 = v_RD_3686_out0;
assign v_RD_3204_out0 = v_RD_3687_out0;
assign v_RD_3208_out0 = v_RD_3689_out0;
assign v_RD_3210_out0 = v_RD_3690_out0;
assign v_RD_3218_out0 = v_RD_3694_out0;
assign v_RD_3220_out0 = v_RD_3695_out0;
assign v_RD_3225_out0 = v_RD_3697_out0;
assign v_RD_3229_out0 = v_RD_3699_out0;
assign v_RD_3231_out0 = v_RD_3700_out0;
assign v_RD_3233_out0 = v_RD_3701_out0;
assign v_RD_3235_out0 = v_RD_3702_out0;
assign v_RD_3239_out0 = v_RD_3704_out0;
assign v_RD_3241_out0 = v_RD_3705_out0;
assign v_RD_3249_out0 = v_RD_3709_out0;
assign v_RD_3251_out0 = v_RD_3710_out0;
assign v_RD_3256_out0 = v_RD_3712_out0;
assign v_RD_3260_out0 = v_RD_3714_out0;
assign v_RD_3262_out0 = v_RD_3715_out0;
assign v_RD_3264_out0 = v_RD_3716_out0;
assign v_RD_3266_out0 = v_RD_3717_out0;
assign v_RD_3270_out0 = v_RD_3719_out0;
assign v_RD_3272_out0 = v_RD_3720_out0;
assign v_RD_3280_out0 = v_RD_3724_out0;
assign v_RD_3282_out0 = v_RD_3725_out0;
assign v_RD_3287_out0 = v_RD_3727_out0;
assign v_RD_3291_out0 = v_RD_3729_out0;
assign v_RD_3293_out0 = v_RD_3730_out0;
assign v_RD_3295_out0 = v_RD_3731_out0;
assign v_RD_3297_out0 = v_RD_3732_out0;
assign v_RD_3301_out0 = v_RD_3734_out0;
assign v_RD_3303_out0 = v_RD_3735_out0;
assign v_RD_3311_out0 = v_RD_3739_out0;
assign v_RD_3313_out0 = v_RD_3740_out0;
assign v_RD_3318_out0 = v_RD_3742_out0;
assign v_RD_3322_out0 = v_RD_3744_out0;
assign v_RD_3324_out0 = v_RD_3745_out0;
assign v_RD_3326_out0 = v_RD_3746_out0;
assign v_RD_3328_out0 = v_RD_3747_out0;
assign v_RD_3332_out0 = v_RD_3749_out0;
assign v_RD_3334_out0 = v_RD_3750_out0;
assign v_RD_3527_out0 = v_G12_6520_out0;
assign v_RD_3528_out0 = v_G14_6735_out0;
assign v_RD_3529_out0 = v_G15_68_out0;
assign v_RD_3532_out0 = v_G13_6577_out0;
assign v_RD_3534_out0 = v_G10_3424_out0;
assign v_RD_3539_out0 = v_G11_315_out0;
assign v_RD_3571_out0 = v_G12_6523_out0;
assign v_RD_3572_out0 = v_G14_6738_out0;
assign v_RD_3573_out0 = v_G15_71_out0;
assign v_RD_3576_out0 = v_G13_6580_out0;
assign v_RD_3578_out0 = v_G10_3427_out0;
assign v_RD_3583_out0 = v_G11_318_out0;
assign v_RD_3601_out0 = v_G12_6525_out0;
assign v_RD_3602_out0 = v_G14_6740_out0;
assign v_RD_3603_out0 = v_G15_73_out0;
assign v_RD_3606_out0 = v_G13_6582_out0;
assign v_RD_3608_out0 = v_G10_3429_out0;
assign v_RD_3613_out0 = v_G11_320_out0;
assign v_RD_3616_out0 = v_G12_6526_out0;
assign v_RD_3617_out0 = v_G14_6741_out0;
assign v_RD_3618_out0 = v_G15_74_out0;
assign v_RD_3621_out0 = v_G13_6583_out0;
assign v_RD_3623_out0 = v_G10_3430_out0;
assign v_RD_3628_out0 = v_G11_321_out0;
assign v_RD_3631_out0 = v_G12_6527_out0;
assign v_RD_3632_out0 = v_G14_6742_out0;
assign v_RD_3633_out0 = v_G15_75_out0;
assign v_RD_3636_out0 = v_G13_6584_out0;
assign v_RD_3638_out0 = v_G10_3431_out0;
assign v_RD_3643_out0 = v_G11_322_out0;
assign v_RD_3646_out0 = v_G12_6528_out0;
assign v_RD_3647_out0 = v_G14_6743_out0;
assign v_RD_3648_out0 = v_G15_76_out0;
assign v_RD_3651_out0 = v_G13_6585_out0;
assign v_RD_3653_out0 = v_G10_3432_out0;
assign v_RD_3658_out0 = v_G11_323_out0;
assign v_RD_3661_out0 = v_G12_6529_out0;
assign v_RD_3662_out0 = v_G14_6744_out0;
assign v_RD_3663_out0 = v_G15_77_out0;
assign v_RD_3666_out0 = v_G13_6586_out0;
assign v_RD_3668_out0 = v_G10_3433_out0;
assign v_RD_3673_out0 = v_G11_324_out0;
assign v_RD_3676_out0 = v_G12_6530_out0;
assign v_RD_3677_out0 = v_G14_6745_out0;
assign v_RD_3678_out0 = v_G15_78_out0;
assign v_RD_3681_out0 = v_G13_6587_out0;
assign v_RD_3683_out0 = v_G10_3434_out0;
assign v_RD_3688_out0 = v_G11_325_out0;
assign v_RD_3691_out0 = v_G12_6531_out0;
assign v_RD_3692_out0 = v_G14_6746_out0;
assign v_RD_3693_out0 = v_G15_79_out0;
assign v_RD_3696_out0 = v_G13_6588_out0;
assign v_RD_3698_out0 = v_G10_3435_out0;
assign v_RD_3703_out0 = v_G11_326_out0;
assign v_RD_3706_out0 = v_G12_6532_out0;
assign v_RD_3707_out0 = v_G14_6747_out0;
assign v_RD_3708_out0 = v_G15_80_out0;
assign v_RD_3711_out0 = v_G13_6589_out0;
assign v_RD_3713_out0 = v_G10_3436_out0;
assign v_RD_3718_out0 = v_G11_327_out0;
assign v_RD_3721_out0 = v_G12_6533_out0;
assign v_RD_3722_out0 = v_G14_6748_out0;
assign v_RD_3723_out0 = v_G15_81_out0;
assign v_RD_3726_out0 = v_G13_6590_out0;
assign v_RD_3728_out0 = v_G10_3437_out0;
assign v_RD_3733_out0 = v_G11_328_out0;
assign v_RD_3736_out0 = v_G12_6534_out0;
assign v_RD_3737_out0 = v_G14_6749_out0;
assign v_RD_3738_out0 = v_G15_82_out0;
assign v_RD_3741_out0 = v_G13_6591_out0;
assign v_RD_3743_out0 = v_G10_3438_out0;
assign v_RD_3748_out0 = v_G11_329_out0;
assign v_ADDER_IN_4304_out0 = v__594_out0;
assign v__5094_out0 = { v_C1_5558_out0,v__5437_out0 };
assign v_MUX1_3_out0 = v_LSL_1388_out0 ? v__5094_out0 : v_IN_4348_out0;
assign v__913_out0 = { v__1310_out0,v__2176_out0 };
assign {v_A1_1547_out1,v_A1_1547_out0 } = v_RM_6657_out0 + v_ADDER_IN_4304_out0 + v_U_5155_out0;
assign v__1905_out0 = v_IN1_1067_out0[0:0];
assign v__1905_out1 = v_IN1_1067_out0[10:10];
assign v_RD_2872_out0 = v_RD_3527_out0;
assign v_RD_2874_out0 = v_RD_3528_out0;
assign v_RD_2876_out0 = v_RD_3529_out0;
assign v_RD_2882_out0 = v_RD_3532_out0;
assign v_RD_2887_out0 = v_RD_3534_out0;
assign v_RD_2897_out0 = v_RD_3539_out0;
assign v_RD_2964_out0 = v_RD_3571_out0;
assign v_RD_2966_out0 = v_RD_3572_out0;
assign v_RD_2968_out0 = v_RD_3573_out0;
assign v_RD_2974_out0 = v_RD_3576_out0;
assign v_RD_2979_out0 = v_RD_3578_out0;
assign v_RD_2989_out0 = v_RD_3583_out0;
assign v_RD_3026_out0 = v_RD_3601_out0;
assign v_RD_3028_out0 = v_RD_3602_out0;
assign v_RD_3030_out0 = v_RD_3603_out0;
assign v_RD_3036_out0 = v_RD_3606_out0;
assign v_RD_3041_out0 = v_RD_3608_out0;
assign v_RD_3051_out0 = v_RD_3613_out0;
assign v_RD_3057_out0 = v_RD_3616_out0;
assign v_RD_3059_out0 = v_RD_3617_out0;
assign v_RD_3061_out0 = v_RD_3618_out0;
assign v_RD_3067_out0 = v_RD_3621_out0;
assign v_RD_3072_out0 = v_RD_3623_out0;
assign v_RD_3082_out0 = v_RD_3628_out0;
assign v_RD_3088_out0 = v_RD_3631_out0;
assign v_RD_3090_out0 = v_RD_3632_out0;
assign v_RD_3092_out0 = v_RD_3633_out0;
assign v_RD_3098_out0 = v_RD_3636_out0;
assign v_RD_3103_out0 = v_RD_3638_out0;
assign v_RD_3113_out0 = v_RD_3643_out0;
assign v_RD_3119_out0 = v_RD_3646_out0;
assign v_RD_3121_out0 = v_RD_3647_out0;
assign v_RD_3123_out0 = v_RD_3648_out0;
assign v_RD_3129_out0 = v_RD_3651_out0;
assign v_RD_3134_out0 = v_RD_3653_out0;
assign v_RD_3144_out0 = v_RD_3658_out0;
assign v_RD_3150_out0 = v_RD_3661_out0;
assign v_RD_3152_out0 = v_RD_3662_out0;
assign v_RD_3154_out0 = v_RD_3663_out0;
assign v_RD_3160_out0 = v_RD_3666_out0;
assign v_RD_3165_out0 = v_RD_3668_out0;
assign v_RD_3175_out0 = v_RD_3673_out0;
assign v_RD_3181_out0 = v_RD_3676_out0;
assign v_RD_3183_out0 = v_RD_3677_out0;
assign v_RD_3185_out0 = v_RD_3678_out0;
assign v_RD_3191_out0 = v_RD_3681_out0;
assign v_RD_3196_out0 = v_RD_3683_out0;
assign v_RD_3206_out0 = v_RD_3688_out0;
assign v_RD_3212_out0 = v_RD_3691_out0;
assign v_RD_3214_out0 = v_RD_3692_out0;
assign v_RD_3216_out0 = v_RD_3693_out0;
assign v_RD_3222_out0 = v_RD_3696_out0;
assign v_RD_3227_out0 = v_RD_3698_out0;
assign v_RD_3237_out0 = v_RD_3703_out0;
assign v_RD_3243_out0 = v_RD_3706_out0;
assign v_RD_3245_out0 = v_RD_3707_out0;
assign v_RD_3247_out0 = v_RD_3708_out0;
assign v_RD_3253_out0 = v_RD_3711_out0;
assign v_RD_3258_out0 = v_RD_3713_out0;
assign v_RD_3268_out0 = v_RD_3718_out0;
assign v_RD_3274_out0 = v_RD_3721_out0;
assign v_RD_3276_out0 = v_RD_3722_out0;
assign v_RD_3278_out0 = v_RD_3723_out0;
assign v_RD_3284_out0 = v_RD_3726_out0;
assign v_RD_3289_out0 = v_RD_3728_out0;
assign v_RD_3299_out0 = v_RD_3733_out0;
assign v_RD_3305_out0 = v_RD_3736_out0;
assign v_RD_3307_out0 = v_RD_3737_out0;
assign v_RD_3309_out0 = v_RD_3738_out0;
assign v_RD_3315_out0 = v_RD_3741_out0;
assign v_RD_3320_out0 = v_RD_3743_out0;
assign v_RD_3330_out0 = v_RD_3748_out0;
assign v_NOTUSED_161_out0 = v__1905_out0;
assign v_ANDOUT_305_out0 = v__913_out0;
assign v__2190_out0 = v_MUX1_3_out0[1:0];
assign v__2190_out1 = v_MUX1_3_out0[15:14];
assign v__2242_out0 = { v__1905_out1,v_C1_4338_out0 };
assign v__2865_out0 = v_A1_1547_out0[11:0];
assign v__2865_out1 = v_A1_1547_out0[15:4];
assign v_COUT_5191_out0 = v_A1_1547_out1;
assign v_RMN_6619_out0 = v_A1_1547_out0;
assign v_OUT1_964_out0 = v__2242_out0;
assign v_NOTUSE_1170_out0 = v__2865_out1;
assign v__5367_out0 = v_ANDOUT_305_out0[0:0];
assign v__5367_out1 = v_ANDOUT_305_out0[15:15];
assign v_UNUSED_5533_out0 = v__2190_out0;
assign v__6641_out0 = { v__2190_out1,v_C1_3337_out0 };
assign v_MUX2_6726_out0 = v_G6_6537_out0 ? v__2865_out0 : v__1479_out0;
assign v_CIN_1148_out0 = v__5367_out1;
assign v_MUX2_5334_out0 = v_LSR_6568_out0 ? v__6641_out0 : v_MUX1_3_out0;
assign v_EA_6661_out0 = v_MUX2_6726_out0;
assign v_MUX5_6734_out0 = v_0_1475_out0 ? v_OUT1_964_out0 : v_IN_6733_out0;
assign v__230_out0 = v_CIN_1148_out0[8:8];
assign v__868_out0 = v_CIN_1148_out0[6:6];
assign v_IN_960_out0 = v_MUX2_5334_out0;
assign v__1051_out0 = v_CIN_1148_out0[3:3];
assign v_RAMADDRMUX_1088_out0 = v_EA_6661_out0;
assign v__1221_out0 = v_CIN_1148_out0[0:0];
assign v__1489_out0 = v_CIN_1148_out0[9:9];
assign v__1505_out0 = v_CIN_1148_out0[2:2];
assign v__1531_out0 = v_CIN_1148_out0[7:7];
assign v__1864_out0 = v_CIN_1148_out0[1:1];
assign v__1882_out0 = v_CIN_1148_out0[10:10];
assign v__3341_out0 = v_CIN_1148_out0[11:11];
assign v__3757_out0 = v_CIN_1148_out0[12:12];
assign v__4283_out0 = v_CIN_1148_out0[13:13];
assign v__4316_out0 = v_CIN_1148_out0[14:14];
assign v__5277_out0 = v_CIN_1148_out0[5:5];
assign v_IN1_5410_out0 = v_MUX5_6734_out0;
assign v__6625_out0 = v_CIN_1148_out0[4:4];
assign v_RAMADDRMUX_48_out0 = v_RAMADDRMUX_1088_out0;
assign v__304_out0 = v_IN_960_out0[1:0];
assign v__304_out1 = v_IN_960_out0[15:14];
assign v_RM_1645_out0 = v__3757_out0;
assign v_RM_1646_out0 = v__4316_out0;
assign v_RM_1647_out0 = v__5277_out0;
assign v_RM_1648_out0 = v__6625_out0;
assign v_RM_1649_out0 = v__4283_out0;
assign v_RM_1650_out0 = v__1489_out0;
assign v_RM_1651_out0 = v__1882_out0;
assign v_RM_1652_out0 = v__1864_out0;
assign v_RM_1653_out0 = v__1051_out0;
assign v_RM_1654_out0 = v__868_out0;
assign v_RM_1655_out0 = v__1531_out0;
assign v_RM_1656_out0 = v__3341_out0;
assign v_RM_1657_out0 = v__230_out0;
assign v_RM_1658_out0 = v__1505_out0;
assign v__5324_out0 = v_IN_960_out0[15:15];
assign v_RM_5604_out0 = v__1221_out0;
assign v__6678_out0 = v_IN1_5410_out0[1:0];
assign v__6678_out1 = v_IN1_5410_out0[10:9];
assign v_NOTUSED_217_out0 = v__6678_out0;
assign v_NOTUSED_218_out0 = v__304_out0;
assign v_G1_3832_out0 = ((v_RD_2913_out0 && !v_RM_5604_out0) || (!v_RD_2913_out0) && v_RM_5604_out0);
assign v__5102_out0 = { v__304_out1,v__5324_out0 };
assign v_RAMADDRMUX_5187_out0 = v_RAMADDRMUX_48_out0;
assign v_RM_5594_out0 = v_RM_1645_out0;
assign v_RM_5596_out0 = v_RM_1646_out0;
assign v_RM_5598_out0 = v_RM_1647_out0;
assign v_RM_5600_out0 = v_RM_1648_out0;
assign v_RM_5602_out0 = v_RM_1649_out0;
assign v_RM_5606_out0 = v_RM_1650_out0;
assign v_RM_5608_out0 = v_RM_1651_out0;
assign v_RM_5610_out0 = v_RM_1652_out0;
assign v_RM_5612_out0 = v_RM_1653_out0;
assign v_RM_5614_out0 = v_RM_1654_out0;
assign v_RM_5616_out0 = v_RM_1655_out0;
assign v_RM_5618_out0 = v_RM_1656_out0;
assign v_RM_5620_out0 = v_RM_1657_out0;
assign v_RM_5622_out0 = v_RM_1658_out0;
assign v_G2_6077_out0 = v_RD_2913_out0 && v_RM_5604_out0;
assign v__6778_out0 = { v__6678_out1,v_C1_1562_out0 };
assign v__575_out0 = { v__5102_out0,v__5324_out0 };
assign v_OUT1_1878_out0 = v__6778_out0;
assign v_CARRY_2414_out0 = v_G2_6077_out0;
assign v_RAMADDRESSMUX_3375_out0 = v_RAMADDRMUX_5187_out0;
assign v_G1_3822_out0 = ((v_RD_2903_out0 && !v_RM_5594_out0) || (!v_RD_2903_out0) && v_RM_5594_out0);
assign v_G1_3824_out0 = ((v_RD_2905_out0 && !v_RM_5596_out0) || (!v_RD_2905_out0) && v_RM_5596_out0);
assign v_G1_3826_out0 = ((v_RD_2907_out0 && !v_RM_5598_out0) || (!v_RD_2907_out0) && v_RM_5598_out0);
assign v_G1_3828_out0 = ((v_RD_2909_out0 && !v_RM_5600_out0) || (!v_RD_2909_out0) && v_RM_5600_out0);
assign v_G1_3830_out0 = ((v_RD_2911_out0 && !v_RM_5602_out0) || (!v_RD_2911_out0) && v_RM_5602_out0);
assign v_G1_3834_out0 = ((v_RD_2915_out0 && !v_RM_5606_out0) || (!v_RD_2915_out0) && v_RM_5606_out0);
assign v_G1_3836_out0 = ((v_RD_2917_out0 && !v_RM_5608_out0) || (!v_RD_2917_out0) && v_RM_5608_out0);
assign v_G1_3838_out0 = ((v_RD_2919_out0 && !v_RM_5610_out0) || (!v_RD_2919_out0) && v_RM_5610_out0);
assign v_G1_3840_out0 = ((v_RD_2921_out0 && !v_RM_5612_out0) || (!v_RD_2921_out0) && v_RM_5612_out0);
assign v_G1_3842_out0 = ((v_RD_2923_out0 && !v_RM_5614_out0) || (!v_RD_2923_out0) && v_RM_5614_out0);
assign v_G1_3844_out0 = ((v_RD_2925_out0 && !v_RM_5616_out0) || (!v_RD_2925_out0) && v_RM_5616_out0);
assign v_G1_3846_out0 = ((v_RD_2927_out0 && !v_RM_5618_out0) || (!v_RD_2927_out0) && v_RM_5618_out0);
assign v_G1_3848_out0 = ((v_RD_2929_out0 && !v_RM_5620_out0) || (!v_RD_2929_out0) && v_RM_5620_out0);
assign v_G1_3850_out0 = ((v_RD_2931_out0 && !v_RM_5622_out0) || (!v_RD_2931_out0) && v_RM_5622_out0);
assign v_RAM_ADDRESS_MUX_4332_out0 = v_RAMADDRMUX_5187_out0;
assign v_S_4401_out0 = v_G1_3832_out0;
assign v_G2_6067_out0 = v_RD_2903_out0 && v_RM_5594_out0;
assign v_G2_6069_out0 = v_RD_2905_out0 && v_RM_5596_out0;
assign v_G2_6071_out0 = v_RD_2907_out0 && v_RM_5598_out0;
assign v_G2_6073_out0 = v_RD_2909_out0 && v_RM_5600_out0;
assign v_G2_6075_out0 = v_RD_2911_out0 && v_RM_5602_out0;
assign v_G2_6079_out0 = v_RD_2915_out0 && v_RM_5606_out0;
assign v_G2_6081_out0 = v_RD_2917_out0 && v_RM_5608_out0;
assign v_G2_6083_out0 = v_RD_2919_out0 && v_RM_5610_out0;
assign v_G2_6085_out0 = v_RD_2921_out0 && v_RM_5612_out0;
assign v_G2_6087_out0 = v_RD_2923_out0 && v_RM_5614_out0;
assign v_G2_6089_out0 = v_RD_2925_out0 && v_RM_5616_out0;
assign v_G2_6091_out0 = v_RD_2927_out0 && v_RM_5618_out0;
assign v_G2_6093_out0 = v_RD_2929_out0 && v_RM_5620_out0;
assign v_G2_6095_out0 = v_RD_2931_out0 && v_RM_5622_out0;
assign v_MUX4_271_out0 = v_1_1860_out0 ? v_OUT1_1878_out0 : v_MUX5_6734_out0;
assign v__1186_out0 = v_RAM_ADDRESS_MUX_4332_out0[3:0];
assign v__1186_out1 = v_RAM_ADDRESS_MUX_4332_out0[11:8];
assign v_S_2279_out0 = v_S_4401_out0;
assign v_CARRY_2404_out0 = v_G2_6067_out0;
assign v_CARRY_2406_out0 = v_G2_6069_out0;
assign v_CARRY_2408_out0 = v_G2_6071_out0;
assign v_CARRY_2410_out0 = v_G2_6073_out0;
assign v_CARRY_2412_out0 = v_G2_6075_out0;
assign v_CARRY_2416_out0 = v_G2_6079_out0;
assign v_CARRY_2418_out0 = v_G2_6081_out0;
assign v_CARRY_2420_out0 = v_G2_6083_out0;
assign v_CARRY_2422_out0 = v_G2_6085_out0;
assign v_CARRY_2424_out0 = v_G2_6087_out0;
assign v_CARRY_2426_out0 = v_G2_6089_out0;
assign v_CARRY_2428_out0 = v_G2_6091_out0;
assign v_CARRY_2430_out0 = v_G2_6093_out0;
assign v_CARRY_2432_out0 = v_G2_6095_out0;
assign v_OUT_4355_out0 = v__575_out0;
assign v_S_4391_out0 = v_G1_3822_out0;
assign v_S_4393_out0 = v_G1_3824_out0;
assign v_S_4395_out0 = v_G1_3826_out0;
assign v_S_4397_out0 = v_G1_3828_out0;
assign v_S_4399_out0 = v_G1_3830_out0;
assign v_S_4403_out0 = v_G1_3834_out0;
assign v_S_4405_out0 = v_G1_3836_out0;
assign v_S_4407_out0 = v_G1_3838_out0;
assign v_S_4409_out0 = v_G1_3840_out0;
assign v_S_4411_out0 = v_G1_3842_out0;
assign v_S_4413_out0 = v_G1_3844_out0;
assign v_S_4415_out0 = v_G1_3846_out0;
assign v_S_4417_out0 = v_G1_3848_out0;
assign v_S_4419_out0 = v_G1_3850_out0;
assign v_CIN_4855_out0 = v_CARRY_2414_out0;
assign v_IN1_1391_out0 = v_MUX4_271_out0;
assign v_MUX3_1527_out0 = v_ASR_6755_out0 ? v_OUT_4355_out0 : v_MUX2_5334_out0;
assign v__1570_out0 = { v__5367_out0,v_S_2279_out0 };
assign v_RD_2920_out0 = v_CIN_4855_out0;
assign v_RM_5595_out0 = v_S_4391_out0;
assign v_RM_5597_out0 = v_S_4393_out0;
assign v_RM_5599_out0 = v_S_4395_out0;
assign v_RM_5601_out0 = v_S_4397_out0;
assign v_RM_5603_out0 = v_S_4399_out0;
assign v_RM_5607_out0 = v_S_4403_out0;
assign v_RM_5609_out0 = v_S_4405_out0;
assign v_RM_5611_out0 = v_S_4407_out0;
assign v_RM_5613_out0 = v_S_4409_out0;
assign v_RM_5615_out0 = v_S_4411_out0;
assign v_RM_5617_out0 = v_S_4413_out0;
assign v_RM_5619_out0 = v_S_4415_out0;
assign v_RM_5621_out0 = v_S_4417_out0;
assign v_RM_5623_out0 = v_S_4419_out0;
assign v__6562_out0 = v__1186_out1[3:0];
assign v__6562_out1 = v__1186_out1[7:4];
assign v_RAM_ADD_BYTE0_6592_out0 = v__1186_out0;
assign v_EQ1_1305_out0 = v__6562_out0 == 4'h1;
assign v__2296_out0 = v_IN1_1391_out0[3:0];
assign v__2296_out1 = v_IN1_1391_out0[10:7];
assign v__2352_out0 = v_MUX3_1527_out0[1:0];
assign v__2352_out1 = v_MUX3_1527_out0[15:14];
assign v_EQ9_2363_out0 = v_RAM_ADD_BYTE0_6592_out0 == 4'h2;
assign v_G1_3839_out0 = ((v_RD_2920_out0 && !v_RM_5611_out0) || (!v_RD_2920_out0) && v_RM_5611_out0);
assign v_EQ01_5173_out0 = v_RAM_ADD_BYTE0_6592_out0 == 4'h1;
assign v_EQ8_5315_out0 = v__6562_out1 == 4'h8;
assign v_G2_6084_out0 = v_RD_2920_out0 && v_RM_5611_out0;
assign v__592_out0 = { v__2352_out1,v__2352_out0 };
assign v_BYTE1_comp1_1189_out0 = v_EQ1_1305_out0;
assign v__1450_out0 = { v__2296_out1,v_C1_5082_out0 };
assign v_CARRY_2421_out0 = v_G2_6084_out0;
assign v_BYTE2_COMP8_3781_out0 = v_EQ8_5315_out0;
assign v_S_4408_out0 = v_G1_3839_out0;
assign v_NOTUSED_5186_out0 = v__2296_out0;
assign v_S_619_out0 = v_S_4408_out0;
assign v_OUT1_916_out0 = v__1450_out0;
assign v_MUX2_1162_out0 = v_BYTE1_comp1_1189_out0 ? v_split_214_out1 : v_split_214_out0;
assign v_G2_1579_out0 = v_EQ01_5173_out0 && v_BYTE2_COMP8_3781_out0;
assign v_G1_1971_out0 = v_CARRY_2421_out0 || v_CARRY_2420_out0;
assign v_MUX4_5179_out0 = v_ROR_1598_out0 ? v__592_out0 : v_MUX3_1527_out0;
assign v_G20_5486_out0 = v_BYTE2_COMP8_3781_out0 && v_EQ9_2363_out0;
assign v_MUX3_6570_out0 = v_BYTE1_comp1_1189_out0 ? v__4824_out0 : v__3476_out0;
assign v_COUT_355_out0 = v_G1_1971_out0;
assign v_MUX5_581_out0 = v_EN_5158_out0 ? v_MUX4_5179_out0 : v_IN_4348_out0;
assign v_TRANSMISSION_DATA_1327_out0 = v_MUX2_1162_out0;
assign v_G14_5126_out0 = v_G2_1579_out0 && v_uart_5478_out0;
assign v_G18_5514_out0 = v_G20_5486_out0 && v_uart_5478_out0;
assign v_REGISTER_TRANSMIT_DATA_6031_out0 = v_MUX2_1162_out0;
assign v_MUX3_6560_out0 = v_2_862_out0 ? v_OUT1_916_out0 : v_MUX4_271_out0;
assign v_TRANSMIT_DATA_39_out0 = v_REGISTER_TRANSMIT_DATA_6031_out0;
assign v_TRANSMISSION_DATA_1422_out0 = v_TRANSMISSION_DATA_1327_out0;
assign v_G19_2277_out0 = v_G18_5514_out0 && v_STORE_110_out0;
assign v_CIN_4861_out0 = v_COUT_355_out0;
assign v_OUT_6029_out0 = v_MUX5_581_out0;
assign v_G16_6595_out0 = v_G14_5126_out0 && v_LOAD_4312_out0;
assign v_IN1_6754_out0 = v_MUX3_6560_out0;
assign v_SEL1_119_out0 = v_TRANSMIT_DATA_39_out0[6:6];
assign v_SEL1_571_out0 = v_TRANSMIT_DATA_39_out0[2:2];
assign v_SEL1_589_out0 = v_TRANSMIT_DATA_39_out0[4:4];
assign v_SEL1_1130_out0 = v_TRANSMIT_DATA_39_out0[0:0];
assign v_SEL1_1183_out0 = v_TRANSMIT_DATA_39_out0[5:5];
assign v_IN_1299_out0 = v_OUT_6029_out0;
assign v__1308_out0 = v_IN1_6754_out0[7:0];
assign v__1308_out1 = v_IN1_6754_out0[10:3];
assign v_G21_1405_out0 = v_G19_2277_out0 && v_EXEC1_1481_out0;
assign v_SEL1_2371_out0 = v_TRANSMIT_DATA_39_out0[3:3];
assign v_RD_2932_out0 = v_CIN_4861_out0;
assign v_SEL1_5081_out0 = v_TRANSMIT_DATA_39_out0[1:1];
assign v_RECEIVING_INSTRUCTION_5497_out0 = v_G16_6595_out0;
assign v_SEL1_6622_out0 = v_TRANSMIT_DATA_39_out0[7:7];
assign v_INSTRUCTION_32_out0 = v_G21_1405_out0;
assign v_RX_INST_49_out0 = v_RECEIVING_INSTRUCTION_5497_out0;
assign v_NOTUSED_331_out0 = v__1308_out0;
assign v__1175_out0 = v_IN_1299_out0[11:0];
assign v__1175_out1 = v_IN_1299_out0[15:4];
assign v_G5_2253_out0 = ! v_RECEIVING_INSTRUCTION_5497_out0;
assign v_G1_3851_out0 = ((v_RD_2932_out0 && !v_RM_5623_out0) || (!v_RD_2932_out0) && v_RM_5623_out0);
assign v_MUX1_5484_out0 = v_RECEIVING_INSTRUCTION_5497_out0 ? v_MUX3_6570_out0 : v_RAM_OUT_5519_out0;
assign v_G2_6096_out0 = v_RD_2932_out0 && v_RM_5623_out0;
assign v__6642_out0 = { v__1308_out1,v_C1_5063_out0 };
assign v_IN_6677_out0 = v_IN_1299_out0;
assign v_G7_17_out0 = v_G6_6648_out0 && v_G5_2253_out0;
assign v_TRANSMIT_INSTRUCTION_839_out0 = v_INSTRUCTION_32_out0;
assign v_NOTUSED1_928_out0 = v__1175_out1;
assign v__1307_out0 = { v_C1_3397_out0,v__1175_out0 };
assign v_RX_INSTRUCTION_1586_out0 = v_RX_INST_49_out0;
assign v_OUT1_1601_out0 = v__6642_out0;
assign v_CARRY_2433_out0 = v_G2_6096_out0;
assign v_TX_INSTRUCTION_3442_out0 = v_INSTRUCTION_32_out0;
assign v_S_4420_out0 = v_G1_3851_out0;
assign v_G3_5370_out0 = v_TX_OVERFLOW_1902_out0 && v_INSTRUCTION_32_out0;
assign v_REGISTER_INPUT_6543_out0 = v_MUX1_5484_out0;
assign v_S_625_out0 = v_S_4420_out0;
assign v_transmit_INSTRUCTION_1304_out0 = v_TRANSMIT_INSTRUCTION_839_out0;
assign v_RAMDOUT_1478_out0 = v_REGISTER_INPUT_6543_out0;
assign v_INSTRCUTION_1926_out0 = v_TX_INSTRUCTION_3442_out0;
assign v_G1_1977_out0 = v_CARRY_2433_out0 || v_CARRY_2432_out0;
assign v_MUX1_2364_out0 = v_LSL_1486_out0 ? v__1307_out0 : v_IN_6677_out0;
assign v_MUX1_3504_out0 = v_3_6711_out0 ? v_OUT1_1601_out0 : v_MUX3_6560_out0;
assign v_G8_6721_out0 = v_G9_1046_out0 || v_G7_17_out0;
assign v_RAMDOUT_14_out0 = v_RAMDOUT_1478_out0;
assign v_COUT_361_out0 = v_G1_1977_out0;
assign v_MUX1_1279_out0 = v_transmit_INSTRUCTION_1304_out0 ? v_SEL1_119_out0 : v_FF1_956_out0;
assign v_shifted1_1300_out0 = v_MUX1_3504_out0;
assign v_MUX8_1316_out0 = v_transmit_INSTRUCTION_1304_out0 ? v_C1_5058_out0 : v_FF8_5523_out0;
assign v_MUX4_1568_out0 = v_transmit_INSTRUCTION_1304_out0 ? v_SEL1_2371_out0 : v_FF4_226_out0;
assign v_MUX2_2175_out0 = v_transmit_INSTRUCTION_1304_out0 ? v_SEL1_1183_out0 : v_FF2_1383_out0;
assign v__2237_out0 = v_MUX1_2364_out0[3:0];
assign v__2237_out1 = v_MUX1_2364_out0[15:12];
assign v__2336_out0 = { v_S_619_out0,v_S_625_out0 };
assign v_MUX3_3503_out0 = v_transmit_INSTRUCTION_1304_out0 ? v_SEL1_589_out0 : v_FF3_5435_out0;
assign v_MUX7_5145_out0 = v_transmit_INSTRUCTION_1304_out0 ? v_SEL1_1130_out0 : v_FF7_2334_out0;
assign v_G2_5156_out0 = ! v_transmit_INSTRUCTION_1304_out0;
assign v_MUX6_5401_out0 = v_transmit_INSTRUCTION_1304_out0 ? v_SEL1_5081_out0 : v_FF6_58_out0;
assign v_MUX5_6574_out0 = v_transmit_INSTRUCTION_1304_out0 ? v_SEL1_571_out0 : v_FF5_3484_out0;
assign v_G3_6656_out0 = v_transmit_INSTRUCTION_1304_out0 || v_SHIFHT_ENABLE_6653_out0;
assign v_G10_292_out0 = v_G7_1195_out0 && v_G2_5156_out0;
assign v_RAMDOUT_1177_out0 = v_RAMDOUT_14_out0;
assign v_ENABLE_1292_out0 = v_G3_6656_out0;
assign v__2276_out0 = { v__2237_out1,v_C1_3397_out0 };
assign v_STARTBIT_3421_out0 = v_G2_5156_out0;
assign v_NOTUSED_4829_out0 = v__2237_out0;
assign v_CIN_4856_out0 = v_COUT_361_out0;
assign v_SHIFTED_SIG_6716_out0 = v_shifted1_1300_out0;
assign v_MUX9_85_out0 = v_G10_292_out0 ? v_2_3472_out0 : v_FF9_4333_out0;
assign v_MUX1_849_out0 = v_EXEC1_12_out0 ? v_RMN_6619_out0 : v_RAMDOUT_1177_out0;
assign v_RD_2922_out0 = v_CIN_4856_out0;
assign v_G35_5105_out0 = v_STARTBIT_3421_out0 && v_G36_1529_out0;
assign v_SHIFTED_SIG_5314_out0 = v_SHIFTED_SIG_6716_out0;
assign v_MUX2_6563_out0 = v_LSR_204_out0 ? v__2276_out0 : v_MUX1_2364_out0;
assign v_MUX2_95_out0 = v_SHIFT_WHICH_OP_2181_out0 ? v_RD_SIG11_3498_out0 : v_SHIFTED_SIG_5314_out0;
assign v_ENABLE_985_out0 = v_G35_5105_out0;
assign v_OUTSTREAM_1024_out0 = v_MUX9_85_out0;
assign v_IN_1145_out0 = v_MUX2_6563_out0;
assign v_MUX1_3784_out0 = v_SHIFT_WHICH_OP_2181_out0 ? v_SHIFTED_SIG_5314_out0 : v_OP2_SIG11_2357_out0;
assign v_G1_3841_out0 = ((v_RD_2922_out0 && !v_RM_5613_out0) || (!v_RD_2922_out0) && v_RM_5613_out0);
assign v_REGDIN_5432_out0 = v_MUX1_849_out0;
assign v_G2_6086_out0 = v_RD_2922_out0 && v_RM_5613_out0;
assign v_OUT_13_out0 = v_OUTSTREAM_1024_out0;
assign v_LS_REGIN_1606_out0 = v_REGDIN_5432_out0;
assign v_CARRY_2423_out0 = v_G2_6086_out0;
assign v_RD_SIG_NEW_4310_out0 = v_MUX2_95_out0;
assign v_G18_4331_out0 = !(v_ENABLE_985_out0 || v_Q7_3383_out0);
assign v_S_4410_out0 = v_G1_3841_out0;
assign v__5184_out0 = v_IN_1145_out0[15:15];
assign v_OP2_SIG_NEW_5507_out0 = v_MUX1_3784_out0;
assign v__6554_out0 = v_IN_1145_out0[3:0];
assign v__6554_out1 = v_IN_1145_out0[15:12];
assign v__84_out0 = { v__6554_out1,v__5184_out0 };
assign v_S_620_out0 = v_S_4410_out0;
assign v_TRANSMITER_1BIT_1200_out0 = v_OUT_13_out0;
assign v_G21_1857_out0 = v_G18_4331_out0 || v_G22_5406_out0;
assign v_G1_1972_out0 = v_CARRY_2423_out0 || v_CARRY_2422_out0;
assign v_RD_SIG_NEW_5348_out0 = v_RD_SIG_NEW_4310_out0;
assign v_OP2_SIG_NEW_5520_out0 = v_OP2_SIG_NEW_5507_out0;
assign v_NOTUSED_6540_out0 = v__6554_out0;
assign v_RD_SIG_56_out0 = v_RD_SIG_NEW_5348_out0;
assign v_COUT_356_out0 = v_G1_1972_out0;
assign v__1245_out0 = { v__2336_out0,v_S_620_out0 };
assign v_TRANSMITER_1BIT_1296_out0 = v_TRANSMITER_1BIT_1200_out0;
assign v__5440_out0 = { v__84_out0,v__5184_out0 };
assign v_OP2_SIG_6561_out0 = v_OP2_SIG_NEW_5520_out0;
assign v__1549_out0 = { v_OP2_SIG_6561_out0,v_C4_1264_out0 };
assign v_CIN_4851_out0 = v_COUT_356_out0;
assign v__5528_out0 = { v__5440_out0,v__5184_out0 };
assign v__6546_out0 = { v_RD_SIG_56_out0,v_C4_1264_out0 };
assign v__1363_out0 = { v__5528_out0,v__5184_out0 };
assign v_XOR2_2192_out0 = v__1549_out0 ^ v_C11_2218_out0;
assign v_RD_2910_out0 = v_CIN_4851_out0;
assign v_XOR1_5534_out0 = v__6546_out0 ^ v_C5_1312_out0;
assign v_OUT_224_out0 = v__1363_out0;
assign {v_A5_929_out1,v_A5_929_out0 } = v_C7_912_out0 + v_XOR2_2192_out0 + v_C12_565_out0;
assign v_G1_3829_out0 = ((v_RD_2910_out0 && !v_RM_5601_out0) || (!v_RD_2910_out0) && v_RM_5601_out0);
assign {v_A4_5526_out1,v_A4_5526_out0 } = v_XOR1_5534_out0 + v_C7_912_out0 + v_C6_5086_out0;
assign v_G2_6074_out0 = v_RD_2910_out0 && v_RM_5601_out0;
assign v_MUX2_579_out0 = v_G1_143_out0 ? v_A5_929_out0 : v__1549_out0;
assign v_MUX1_921_out0 = v_RD_SIGN_1173_out0 ? v_A4_5526_out0 : v__6546_out0;
assign v_MUX3_1483_out0 = v_ASR_5199_out0 ? v_OUT_224_out0 : v_MUX2_6563_out0;
assign v_CARRY_2411_out0 = v_G2_6074_out0;
assign v_S_4398_out0 = v_G1_3829_out0;
assign v_NOTUSED4_5182_out0 = v_A4_5526_out1;
assign v_NOTUSED1_5259_out0 = v_A5_929_out1;
assign v_S_615_out0 = v_S_4398_out0;
assign v_G1_1967_out0 = v_CARRY_2411_out0 || v_CARRY_2410_out0;
assign v__2193_out0 = v_MUX3_1483_out0[3:0];
assign v__2193_out1 = v_MUX3_1483_out0[15:12];
assign {v_A6_5152_out1,v_A6_5152_out0 } = v_MUX1_921_out0 + v_MUX2_579_out0 + v_C3_2314_out0;
assign v__86_out0 = { v__2193_out1,v__2193_out0 };
assign v_COUT_351_out0 = v_G1_1967_out0;
assign v_SEL1_1125_out0 = v_A6_5152_out0[15:15];
assign v__3453_out0 = { v__1245_out0,v_S_615_out0 };
assign v_NOTUSED_5331_out0 = v_A6_5152_out1;
assign v_XOR3_6702_out0 = v_A6_5152_out0 ^ v_C15_847_out0;
assign v_SIGN_ANS_963_out0 = v_SEL1_1125_out0;
assign v_MUX4_1087_out0 = v_ROR_267_out0 ? v__86_out0 : v_MUX3_1483_out0;
assign v_CIN_4850_out0 = v_COUT_351_out0;
assign {v_A8_5490_out1,v_A8_5490_out0 } = v_XOR3_6702_out0 + v_C13_1065_out0 + v_C14_822_out0;
assign v_NOTUSED2_2839_out0 = v_A8_5490_out1;
assign v_RD_2908_out0 = v_CIN_4850_out0;
assign v_SIGN_ANS_4257_out0 = v_SIGN_ANS_963_out0;
assign v_MUX3_4267_out0 = v_SEL1_1125_out0 ? v_A8_5490_out0 : v_A6_5152_out0;
assign v_MUX5_5220_out0 = v_EN_6500_out0 ? v_MUX4_1087_out0 : v_IN_6677_out0;
assign v_OUT_1146_out0 = v_MUX5_5220_out0;
assign v_SIGN_ANS_2180_out0 = v_SIGN_ANS_4257_out0;
assign v_G1_3827_out0 = ((v_RD_2908_out0 && !v_RM_5599_out0) || (!v_RD_2908_out0) && v_RM_5599_out0);
assign v_SEL8_5260_out0 = v_MUX3_4267_out0[11:0];
assign v_G2_6072_out0 = v_RD_2908_out0 && v_RM_5599_out0;
assign v_IN_96_out0 = v_OUT_1146_out0;
assign v_CARRY_2409_out0 = v_G2_6072_out0;
assign v_S_4396_out0 = v_G1_3827_out0;
assign v_SIGN_ANS_5080_out0 = v_SIGN_ANS_2180_out0;
assign v_IN_332_out0 = v_IN_96_out0;
assign v_S_614_out0 = v_S_4396_out0;
assign v__1524_out0 = v_IN_96_out0[7:0];
assign v__1524_out1 = v_IN_96_out0[15:8];
assign v_G1_1966_out0 = v_CARRY_2409_out0 || v_CARRY_2408_out0;
assign v_NOTUSED2_23_out0 = v__1524_out1;
assign v_COUT_350_out0 = v_G1_1966_out0;
assign v__2299_out0 = { v_C1_6623_out0,v__1524_out0 };
assign v__6663_out0 = { v__3453_out0,v_S_614_out0 };
assign v_CIN_4857_out0 = v_COUT_350_out0;
assign v_MUX1_5143_out0 = v_LSL_909_out0 ? v__2299_out0 : v_IN_332_out0;
assign v_RD_2924_out0 = v_CIN_4857_out0;
assign v__4270_out0 = v_MUX1_5143_out0[7:0];
assign v__4270_out1 = v_MUX1_5143_out0[15:8];
assign v_G1_3843_out0 = ((v_RD_2924_out0 && !v_RM_5615_out0) || (!v_RD_2924_out0) && v_RM_5615_out0);
assign v__5170_out0 = { v__4270_out1,v_C1_6623_out0 };
assign v_NOTUSED_5198_out0 = v__4270_out0;
assign v_G2_6088_out0 = v_RD_2924_out0 && v_RM_5615_out0;
assign v_MUX2_1140_out0 = v_LSR_576_out0 ? v__5170_out0 : v_MUX1_5143_out0;
assign v_CARRY_2425_out0 = v_G2_6088_out0;
assign v_S_4412_out0 = v_G1_3843_out0;
assign v_S_621_out0 = v_S_4412_out0;
assign v_G1_1973_out0 = v_CARRY_2425_out0 || v_CARRY_2424_out0;
assign v_IN_2840_out0 = v_MUX2_1140_out0;
assign v_COUT_357_out0 = v_G1_1973_out0;
assign v__1259_out0 = v_IN_2840_out0[7:0];
assign v__1259_out1 = v_IN_2840_out0[15:8];
assign v__1588_out0 = v_IN_2840_out0[15:15];
assign v__1611_out0 = { v__6663_out0,v_S_621_out0 };
assign v_NOTUSED_35_out0 = v__1259_out0;
assign v__3785_out0 = { v__1259_out1,v__1588_out0 };
assign v_CIN_4858_out0 = v_COUT_357_out0;
assign v_RD_2926_out0 = v_CIN_4858_out0;
assign v__5316_out0 = { v__3785_out0,v__1588_out0 };
assign v_G1_3845_out0 = ((v_RD_2926_out0 && !v_RM_5617_out0) || (!v_RD_2926_out0) && v_RM_5617_out0);
assign v_G2_6090_out0 = v_RD_2926_out0 && v_RM_5617_out0;
assign v__6559_out0 = { v__5316_out0,v__1588_out0 };
assign v__55_out0 = { v__6559_out0,v__1588_out0 };
assign v_CARRY_2427_out0 = v_G2_6090_out0;
assign v_S_4414_out0 = v_G1_3845_out0;
assign v_S_622_out0 = v_S_4414_out0;
assign v_G1_1974_out0 = v_CARRY_2427_out0 || v_CARRY_2426_out0;
assign v__2867_out0 = { v__55_out0,v__1588_out0 };
assign v__264_out0 = { v__2867_out0,v__1588_out0 };
assign v_COUT_358_out0 = v_G1_1974_out0;
assign v__3508_out0 = { v__1611_out0,v_S_622_out0 };
assign v__1084_out0 = { v__264_out0,v__1588_out0 };
assign v_CIN_4860_out0 = v_COUT_358_out0;
assign v_RD_2930_out0 = v_CIN_4860_out0;
assign v__3494_out0 = { v__1084_out0,v__1588_out0 };
assign v_OUT_1394_out0 = v__3494_out0;
assign v_G1_3849_out0 = ((v_RD_2930_out0 && !v_RM_5621_out0) || (!v_RD_2930_out0) && v_RM_5621_out0);
assign v_G2_6094_out0 = v_RD_2930_out0 && v_RM_5621_out0;
assign v_CARRY_2431_out0 = v_G2_6094_out0;
assign v_MUX3_3371_out0 = v_ASR_5107_out0 ? v_OUT_1394_out0 : v_MUX2_1140_out0;
assign v_S_4418_out0 = v_G1_3849_out0;
assign v_S_624_out0 = v_S_4418_out0;
assign v_G1_1976_out0 = v_CARRY_2431_out0 || v_CARRY_2430_out0;
assign v__5480_out0 = v_MUX3_3371_out0[7:0];
assign v__5480_out1 = v_MUX3_3371_out0[15:8];
assign v_COUT_360_out0 = v_G1_1976_out0;
assign v__2319_out0 = { v__3508_out0,v_S_624_out0 };
assign v__3374_out0 = { v__5480_out1,v__5480_out0 };
assign v_CIN_4853_out0 = v_COUT_360_out0;
assign v_MUX4_6651_out0 = v_ROR_140_out0 ? v__3374_out0 : v_MUX3_3371_out0;
assign v_MUX5_1607_out0 = v_EN_1190_out0 ? v_MUX4_6651_out0 : v_IN_332_out0;
assign v_RD_2916_out0 = v_CIN_4853_out0;
assign v_G1_3835_out0 = ((v_RD_2916_out0 && !v_RM_5607_out0) || (!v_RD_2916_out0) && v_RM_5607_out0);
assign v_OUT_5062_out0 = v_MUX5_1607_out0;
assign v_G2_6080_out0 = v_RD_2916_out0 && v_RM_5607_out0;
assign v_OP2_1397_out0 = v_OUT_5062_out0;
assign v_CARRY_2417_out0 = v_G2_6080_out0;
assign v_S_4404_out0 = v_G1_3835_out0;
assign v_S_617_out0 = v_S_4404_out0;
assign v_G1_1969_out0 = v_CARRY_2417_out0 || v_CARRY_2416_out0;
assign v_OP2_5489_out0 = v_OP2_1397_out0;
assign v_COUT_353_out0 = v_G1_1969_out0;
assign v_OP2_1921_out0 = v_OP2_5489_out0;
assign v__3401_out0 = { v__2319_out0,v_S_617_out0 };
assign v_OP2_1132_out0 = v_OP2_1921_out0;
assign v_CIN_4854_out0 = v_COUT_353_out0;
assign v_RD_2918_out0 = v_CIN_4854_out0;
assign v_OP2_5292_out0 = v_OP2_1132_out0;
assign v_MUX5_1265_out0 = v_MOV_99_out0 ? v_OP2_5292_out0 : v_OP1_1005_out0;
assign v_B_1629_out0 = v_OP2_5292_out0;
assign v_G1_3837_out0 = ((v_RD_2918_out0 && !v_RM_5609_out0) || (!v_RD_2918_out0) && v_RM_5609_out0);
assign v_A_5537_out0 = v_OP2_5292_out0;
assign v_G2_6082_out0 = v_RD_2918_out0 && v_RM_5609_out0;
assign v__40_out0 = v_A_5537_out0[3:3];
assign v__97_out0 = v_A_5537_out0[15:15];
assign v__100_out0 = v_B_1629_out0[7:7];
assign v__159_out0 = v_A_5537_out0[0:0];
assign v__163_out0 = v_A_5537_out0[9:9];
assign v__844_out0 = v_B_1629_out0[5:5];
assign v__931_out0 = v_B_1629_out0[9:9];
assign v__1022_out0 = v_A_5537_out0[13:13];
assign v__1179_out0 = v_A_5537_out0[6:6];
assign v__1199_out0 = v_B_1629_out0[2:2];
assign v__1436_out0 = v_B_1629_out0[10:10];
assign v__1521_out0 = v_A_5537_out0[14:14];
assign v__1576_out0 = v_B_1629_out0[11:11];
assign v__1596_out0 = v_A_5537_out0[2:2];
assign v__2251_out0 = v_B_1629_out0[3:3];
assign v__2350_out0 = v_B_1629_out0[4:4];
assign v__2351_out0 = v_B_1629_out0[14:14];
assign v__2359_out0 = v_B_1629_out0[6:6];
assign v_CARRY_2419_out0 = v_G2_6082_out0;
assign v__3471_out0 = v_B_1629_out0[0:0];
assign v__4305_out0 = v_A_5537_out0[8:8];
assign v__4343_out0 = v_A_5537_out0[7:7];
assign v__4345_out0 = v_B_1629_out0[15:15];
assign v_S_4406_out0 = v_G1_3837_out0;
assign v__5111_out0 = v_A_5537_out0[5:5];
assign v__5115_out0 = v_A_5537_out0[1:1];
assign v__5185_out0 = v_B_1629_out0[13:13];
assign v__5264_out0 = v_A_5537_out0[4:4];
assign v__5304_out0 = v_A_5537_out0[12:12];
assign v__5343_out0 = v_A_5537_out0[10:10];
assign v__5518_out0 = v_B_1629_out0[12:12];
assign v__6535_out0 = v_B_1629_out0[1:1];
assign v__6597_out0 = v_B_1629_out0[8:8];
assign v__6679_out0 = v_A_5537_out0[11:11];
assign v_G3_103_out0 = ((v__1596_out0 && !v_SUB_2255_out0) || (!v__1596_out0) && v_SUB_2255_out0);
assign v_G8_270_out0 = v__6594_out0 && v__100_out0;
assign v_G14_299_out0 = v__2301_out0 && v__5185_out0;
assign v_G13_311_out0 = v__1402_out0 && v__5518_out0;
assign v_G8_595_out0 = ((v__4343_out0 && !v_SUB_2255_out0) || (!v__4343_out0) && v_SUB_2255_out0);
assign v_S_618_out0 = v_S_4406_out0;
assign v_G2_885_out0 = v__6660_out0 && v__6535_out0;
assign v_G15_886_out0 = ((v__1521_out0 && !v_SUB_2255_out0) || (!v__1521_out0) && v_SUB_2255_out0);
assign v_G1_920_out0 = v__927_out0 && v__3471_out0;
assign v_G10_1288_out0 = v__6715_out0 && v__931_out0;
assign v_G4_1351_out0 = v__1404_out0 && v__2251_out0;
assign v_G7_1356_out0 = ((v__1179_out0 && !v_SUB_2255_out0) || (!v__1179_out0) && v_SUB_2255_out0);
assign v_G5_1359_out0 = v__1_out0 && v__2350_out0;
assign v_G9_1411_out0 = v__1581_out0 && v__6597_out0;
assign v_G11_1434_out0 = v__2245_out0 && v__1436_out0;
assign v_G12_1626_out0 = ((v__6679_out0 && !v_SUB_2255_out0) || (!v__6679_out0) && v_SUB_2255_out0);
assign v_G1_1970_out0 = v_CARRY_2419_out0 || v_CARRY_2418_out0;
assign v_G14_2215_out0 = ((v__1022_out0 && !v_SUB_2255_out0) || (!v__1022_out0) && v_SUB_2255_out0);
assign v_G15_2275_out0 = v__4354_out0 && v__2351_out0;
assign v_G13_2297_out0 = ((v__5304_out0 && !v_SUB_2255_out0) || (!v__5304_out0) && v_SUB_2255_out0);
assign v_G2_3449_out0 = ((v__5115_out0 && !v_SUB_2255_out0) || (!v__5115_out0) && v_SUB_2255_out0);
assign v_G3_3480_out0 = v__1049_out0 && v__1199_out0;
assign v_G7_4261_out0 = v__5488_out0 && v__2359_out0;
assign v_G6_4347_out0 = v__832_out0 && v__844_out0;
assign v_G5_5200_out0 = ((v__5264_out0 && !v_SUB_2255_out0) || (!v__5264_out0) && v_SUB_2255_out0);
assign v_G12_5262_out0 = v__854_out0 && v__1576_out0;
assign v_G16_5366_out0 = v__1348_out0 && v__4345_out0;
assign v_G4_5412_out0 = ((v__40_out0 && !v_SUB_2255_out0) || (!v__40_out0) && v_SUB_2255_out0);
assign v_G16_5430_out0 = ((v__97_out0 && !v_SUB_2255_out0) || (!v__97_out0) && v_SUB_2255_out0);
assign v_G10_6517_out0 = ((v__163_out0 && !v_SUB_2255_out0) || (!v__163_out0) && v_SUB_2255_out0);
assign v_G9_6551_out0 = ((v__4305_out0 && !v_SUB_2255_out0) || (!v__4305_out0) && v_SUB_2255_out0);
assign v_G11_6572_out0 = ((v__5343_out0 && !v_SUB_2255_out0) || (!v__5343_out0) && v_SUB_2255_out0);
assign v_G6_6718_out0 = ((v__5111_out0 && !v_SUB_2255_out0) || (!v__5111_out0) && v_SUB_2255_out0);
assign v_G1_6776_out0 = ((v__159_out0 && !v_SUB_2255_out0) || (!v__159_out0) && v_SUB_2255_out0);
assign v__189_out0 = { v_G5_1359_out0,v_G6_4347_out0 };
assign v__194_out0 = { v_G9_1411_out0,v_G10_1288_out0 };
assign v_COUT_354_out0 = v_G1_1970_out0;
assign v__954_out0 = { v_G1_6776_out0,v_G2_3449_out0 };
assign v__1438_out0 = { v_G15_2275_out0,v_G16_5366_out0 };
assign v__1567_out0 = { v_G1_920_out0,v_G2_885_out0 };
assign v__1595_out0 = { v_G3_3480_out0,v_G4_1351_out0 };
assign v__2845_out0 = { v__3401_out0,v_S_618_out0 };
assign v__3502_out0 = { v_G13_311_out0,v_G14_299_out0 };
assign v__6539_out0 = { v_G11_1434_out0,v_G12_5262_out0 };
assign v__6784_out0 = { v_G7_4261_out0,v_G8_270_out0 };
assign v__60_out0 = { v__189_out0,v__6784_out0 };
assign v__220_out0 = { v__3502_out0,v__1438_out0 };
assign v__1144_out0 = { v__194_out0,v__6539_out0 };
assign v__4831_out0 = { v__954_out0,v_G3_103_out0 };
assign v_CIN_4859_out0 = v_COUT_354_out0;
assign v__5110_out0 = { v__1567_out0,v__1595_out0 };
assign v__1311_out0 = { v__5110_out0,v__60_out0 };
assign v__2177_out0 = { v__1144_out0,v__220_out0 };
assign v_RD_2928_out0 = v_CIN_4859_out0;
assign v__4276_out0 = { v__4831_out0,v_G4_5412_out0 };
assign v__914_out0 = { v__1311_out0,v__2177_out0 };
assign v__1583_out0 = { v__4276_out0,v_G5_5200_out0 };
assign v_G1_3847_out0 = ((v_RD_2928_out0 && !v_RM_5619_out0) || (!v_RD_2928_out0) && v_RM_5619_out0);
assign v_G2_6092_out0 = v_RD_2928_out0 && v_RM_5619_out0;
assign v_ANDOUT_306_out0 = v__914_out0;
assign v_CARRY_2429_out0 = v_G2_6092_out0;
assign v_S_4416_out0 = v_G1_3847_out0;
assign v__5078_out0 = { v__1583_out0,v_G6_6718_out0 };
assign v__62_out0 = { v__5078_out0,v_G7_1356_out0 };
assign v_S_623_out0 = v_S_4416_out0;
assign v_G1_1975_out0 = v_CARRY_2429_out0 || v_CARRY_2428_out0;
assign v_COUT_359_out0 = v_G1_1975_out0;
assign v__989_out0 = { v__2845_out0,v_S_623_out0 };
assign v__6793_out0 = { v__62_out0,v_G8_595_out0 };
assign v__227_out0 = { v__6793_out0,v_G9_6551_out0 };
assign v_CIN_4848_out0 = v_COUT_359_out0;
assign v__206_out0 = { v__227_out0,v_G10_6517_out0 };
assign v_RD_2904_out0 = v_CIN_4848_out0;
assign v__1384_out0 = { v__206_out0,v_G11_6572_out0 };
assign v_G1_3823_out0 = ((v_RD_2904_out0 && !v_RM_5595_out0) || (!v_RD_2904_out0) && v_RM_5595_out0);
assign v_G2_6068_out0 = v_RD_2904_out0 && v_RM_5595_out0;
assign v_CARRY_2405_out0 = v_G2_6068_out0;
assign v_S_4392_out0 = v_G1_3823_out0;
assign v__5482_out0 = { v__1384_out0,v_G12_1626_out0 };
assign v_S_612_out0 = v_S_4392_out0;
assign v__1557_out0 = { v__5482_out0,v_G13_2297_out0 };
assign v_G1_1964_out0 = v_CARRY_2405_out0 || v_CARRY_2404_out0;
assign v__89_out0 = { v__1557_out0,v_G14_2215_out0 };
assign v_COUT_348_out0 = v_G1_1964_out0;
assign v__1365_out0 = { v__989_out0,v_S_612_out0 };
assign v_CIN_4852_out0 = v_COUT_348_out0;
assign v__5149_out0 = { v__89_out0,v_G15_886_out0 };
assign v__593_out0 = { v__5149_out0,v_G16_5430_out0 };
assign v_RD_2912_out0 = v_CIN_4852_out0;
assign v_G1_3831_out0 = ((v_RD_2912_out0 && !v_RM_5603_out0) || (!v_RD_2912_out0) && v_RM_5603_out0);
assign v_ADDER_IN_4303_out0 = v__593_out0;
assign v_G2_6076_out0 = v_RD_2912_out0 && v_RM_5603_out0;
assign {v_A1_1879_out1,v_A1_1879_out0 } = v_OP1_1005_out0 + v_ADDER_IN_4303_out0 + v_G10_67_out0;
assign v_CARRY_2413_out0 = v_G2_6076_out0;
assign v_S_4400_out0 = v_G1_3831_out0;
assign v_S_616_out0 = v_S_4400_out0;
assign v_COUT_1898_out0 = v_A1_1879_out1;
assign v_G1_1968_out0 = v_CARRY_2413_out0 || v_CARRY_2412_out0;
assign v_SUM1_6516_out0 = v_A1_1879_out0;
assign v_COUT_352_out0 = v_G1_1968_out0;
assign v__892_out0 = { v__1365_out0,v_S_616_out0 };
assign v_MUX3_1004_out0 = v_G7_87_out0 ? v_SUM1_6516_out0 : v_MUX5_1265_out0;
assign v_MUX2_588_out0 = v_G9_199_out0 ? v_ANDOUT_306_out0 : v_MUX3_1004_out0;
assign v_CIN_4849_out0 = v_COUT_352_out0;
assign v_RD_2906_out0 = v_CIN_4849_out0;
assign v_ALUOUT_5181_out0 = v_MUX2_588_out0;
assign v_G1_3825_out0 = ((v_RD_2906_out0 && !v_RM_5597_out0) || (!v_RD_2906_out0) && v_RM_5597_out0);
assign v_ALUOUT_4357_out0 = v_ALUOUT_5181_out0;
assign v_G2_6070_out0 = v_RD_2906_out0 && v_RM_5597_out0;
assign v_ALUOUT_2249_out0 = v_ALUOUT_4357_out0;
assign v_CARRY_2407_out0 = v_G2_6070_out0;
assign v_S_4394_out0 = v_G1_3825_out0;
assign v_S_613_out0 = v_S_4394_out0;
assign v_G1_1965_out0 = v_CARRY_2407_out0 || v_CARRY_2406_out0;
assign v_ALUOUT_5439_out0 = v_ALUOUT_2249_out0;
assign v_COUT_349_out0 = v_G1_1965_out0;
assign v_ALUOUT_2195_out0 = v_ALUOUT_5439_out0;
assign v__2221_out0 = { v__892_out0,v_S_613_out0 };
assign v_EQ3_5434_out0 = v_ALUOUT_2195_out0 == 16'h0;
assign v__5559_out0 = v_ALUOUT_2195_out0[14:0];
assign v__5559_out1 = v_ALUOUT_2195_out0[15:1];
assign v_RM_5605_out0 = v_COUT_349_out0;
assign v_EQ_52_out0 = v_EQ3_5434_out0;
assign v_REST_83_out0 = v__5559_out0;
assign v_MI_1273_out0 = v__5559_out1;
assign v_G1_3833_out0 = ((v_RD_2914_out0 && !v_RM_5605_out0) || (!v_RD_2914_out0) && v_RM_5605_out0);
assign v_G2_6078_out0 = v_RD_2914_out0 && v_RM_5605_out0;
assign v_MI_274_out0 = v_MI_1273_out0;
assign v_EQ_1263_out0 = v_EQ_52_out0;
assign v_CARRY_2415_out0 = v_G2_6078_out0;
assign v_S_4402_out0 = v_G1_3833_out0;
assign v_EQ_1862_out0 = v_EQ_1263_out0;
assign v__5244_out0 = { v__2221_out0,v_S_4402_out0 };
assign v_MI_5330_out0 = v_MI_274_out0;
assign v_JMIN_1298_out0 = v_MI_5330_out0;
assign v_JEQZ_5174_out0 = v_EQ_1862_out0;
assign v__5387_out0 = { v__5244_out0,v_CARRY_2415_out0 };
assign v_JMIN_590_out0 = v_JMIN_1298_out0;
assign v_JEQZ_1455_out0 = v_JEQZ_5174_out0;
assign v_COUT_5372_out0 = v__5387_out0;
assign v_CIN_1149_out0 = v_COUT_5372_out0;
assign v_G4_2365_out0 = v_JEQZ_1455_out0 && v_JEQ_4334_out0;
assign v_G5_5183_out0 = v_JMIN_590_out0 && v_JMI_1565_out0;
assign v__231_out0 = v_CIN_1149_out0[8:8];
assign v__869_out0 = v_CIN_1149_out0[6:6];
assign v__1052_out0 = v_CIN_1149_out0[3:3];
assign v__1071_out0 = v_CIN_1149_out0[15:15];
assign v__1222_out0 = v_CIN_1149_out0[0:0];
assign v__1490_out0 = v_CIN_1149_out0[9:9];
assign v__1506_out0 = v_CIN_1149_out0[2:2];
assign v__1532_out0 = v_CIN_1149_out0[7:7];
assign v__1865_out0 = v_CIN_1149_out0[1:1];
assign v__1883_out0 = v_CIN_1149_out0[10:10];
assign v__3342_out0 = v_CIN_1149_out0[11:11];
assign v__3758_out0 = v_CIN_1149_out0[12:12];
assign v__4284_out0 = v_CIN_1149_out0[13:13];
assign v__4317_out0 = v_CIN_1149_out0[14:14];
assign v__5278_out0 = v_CIN_1149_out0[5:5];
assign v__6626_out0 = v_CIN_1149_out0[4:4];
assign v_G2_6723_out0 = v_JMP_268_out0 || v_G5_5183_out0;
assign v_RM_1659_out0 = v__3758_out0;
assign v_RM_1660_out0 = v__4317_out0;
assign v_RM_1662_out0 = v__5278_out0;
assign v_RM_1663_out0 = v__6626_out0;
assign v_RM_1664_out0 = v__4284_out0;
assign v_RM_1665_out0 = v__1490_out0;
assign v_RM_1666_out0 = v__1883_out0;
assign v_RM_1667_out0 = v__1865_out0;
assign v_RM_1668_out0 = v__1052_out0;
assign v_RM_1669_out0 = v__869_out0;
assign v_RM_1670_out0 = v__1532_out0;
assign v_RM_1671_out0 = v__3342_out0;
assign v_RM_1672_out0 = v__231_out0;
assign v_RM_1673_out0 = v__1506_out0;
assign v_G3_1858_out0 = v_G2_6723_out0 || v_G4_2365_out0;
assign v_CIN_4864_out0 = v__1071_out0;
assign v_RM_5636_out0 = v__1222_out0;
assign v_JUMP_1066_out0 = v_G3_1858_out0;
assign v_RD_2938_out0 = v_CIN_4864_out0;
assign v_G1_3864_out0 = ((v_RD_2945_out0 && !v_RM_5636_out0) || (!v_RD_2945_out0) && v_RM_5636_out0);
assign v_RM_5624_out0 = v_RM_1659_out0;
assign v_RM_5626_out0 = v_RM_1660_out0;
assign v_RM_5630_out0 = v_RM_1662_out0;
assign v_RM_5632_out0 = v_RM_1663_out0;
assign v_RM_5634_out0 = v_RM_1664_out0;
assign v_RM_5637_out0 = v_RM_1665_out0;
assign v_RM_5639_out0 = v_RM_1666_out0;
assign v_RM_5641_out0 = v_RM_1667_out0;
assign v_RM_5643_out0 = v_RM_1668_out0;
assign v_RM_5645_out0 = v_RM_1669_out0;
assign v_RM_5647_out0 = v_RM_1670_out0;
assign v_RM_5649_out0 = v_RM_1671_out0;
assign v_RM_5651_out0 = v_RM_1672_out0;
assign v_RM_5653_out0 = v_RM_1673_out0;
assign v_G2_6109_out0 = v_RD_2945_out0 && v_RM_5636_out0;
assign v_G14_578_out0 = v_G15_906_out0 && v_JUMP_1066_out0;
assign v_CARRY_2446_out0 = v_G2_6109_out0;
assign v_G1_3852_out0 = ((v_RD_2933_out0 && !v_RM_5624_out0) || (!v_RD_2933_out0) && v_RM_5624_out0);
assign v_G1_3854_out0 = ((v_RD_2935_out0 && !v_RM_5626_out0) || (!v_RD_2935_out0) && v_RM_5626_out0);
assign v_G1_3858_out0 = ((v_RD_2939_out0 && !v_RM_5630_out0) || (!v_RD_2939_out0) && v_RM_5630_out0);
assign v_G1_3860_out0 = ((v_RD_2941_out0 && !v_RM_5632_out0) || (!v_RD_2941_out0) && v_RM_5632_out0);
assign v_G1_3862_out0 = ((v_RD_2943_out0 && !v_RM_5634_out0) || (!v_RD_2943_out0) && v_RM_5634_out0);
assign v_G1_3865_out0 = ((v_RD_2946_out0 && !v_RM_5637_out0) || (!v_RD_2946_out0) && v_RM_5637_out0);
assign v_G1_3867_out0 = ((v_RD_2948_out0 && !v_RM_5639_out0) || (!v_RD_2948_out0) && v_RM_5639_out0);
assign v_G1_3869_out0 = ((v_RD_2950_out0 && !v_RM_5641_out0) || (!v_RD_2950_out0) && v_RM_5641_out0);
assign v_G1_3871_out0 = ((v_RD_2952_out0 && !v_RM_5643_out0) || (!v_RD_2952_out0) && v_RM_5643_out0);
assign v_G1_3873_out0 = ((v_RD_2954_out0 && !v_RM_5645_out0) || (!v_RD_2954_out0) && v_RM_5645_out0);
assign v_G1_3875_out0 = ((v_RD_2956_out0 && !v_RM_5647_out0) || (!v_RD_2956_out0) && v_RM_5647_out0);
assign v_G1_3877_out0 = ((v_RD_2958_out0 && !v_RM_5649_out0) || (!v_RD_2958_out0) && v_RM_5649_out0);
assign v_G1_3879_out0 = ((v_RD_2960_out0 && !v_RM_5651_out0) || (!v_RD_2960_out0) && v_RM_5651_out0);
assign v_G1_3881_out0 = ((v_RD_2962_out0 && !v_RM_5653_out0) || (!v_RD_2962_out0) && v_RM_5653_out0);
assign v_S_4433_out0 = v_G1_3864_out0;
assign v_G2_6097_out0 = v_RD_2933_out0 && v_RM_5624_out0;
assign v_G2_6099_out0 = v_RD_2935_out0 && v_RM_5626_out0;
assign v_G2_6103_out0 = v_RD_2939_out0 && v_RM_5630_out0;
assign v_G2_6105_out0 = v_RD_2941_out0 && v_RM_5632_out0;
assign v_G2_6107_out0 = v_RD_2943_out0 && v_RM_5634_out0;
assign v_G2_6110_out0 = v_RD_2946_out0 && v_RM_5637_out0;
assign v_G2_6112_out0 = v_RD_2948_out0 && v_RM_5639_out0;
assign v_G2_6114_out0 = v_RD_2950_out0 && v_RM_5641_out0;
assign v_G2_6116_out0 = v_RD_2952_out0 && v_RM_5643_out0;
assign v_G2_6118_out0 = v_RD_2954_out0 && v_RM_5645_out0;
assign v_G2_6120_out0 = v_RD_2956_out0 && v_RM_5647_out0;
assign v_G2_6122_out0 = v_RD_2958_out0 && v_RM_5649_out0;
assign v_G2_6124_out0 = v_RD_2960_out0 && v_RM_5651_out0;
assign v_G2_6126_out0 = v_RD_2962_out0 && v_RM_5653_out0;
assign v_S_2280_out0 = v_S_4433_out0;
assign v_CARRY_2434_out0 = v_G2_6097_out0;
assign v_CARRY_2436_out0 = v_G2_6099_out0;
assign v_CARRY_2440_out0 = v_G2_6103_out0;
assign v_CARRY_2442_out0 = v_G2_6105_out0;
assign v_CARRY_2444_out0 = v_G2_6107_out0;
assign v_CARRY_2447_out0 = v_G2_6110_out0;
assign v_CARRY_2449_out0 = v_G2_6112_out0;
assign v_CARRY_2451_out0 = v_G2_6114_out0;
assign v_CARRY_2453_out0 = v_G2_6116_out0;
assign v_CARRY_2455_out0 = v_G2_6118_out0;
assign v_CARRY_2457_out0 = v_G2_6120_out0;
assign v_CARRY_2459_out0 = v_G2_6122_out0;
assign v_CARRY_2461_out0 = v_G2_6124_out0;
assign v_CARRY_2463_out0 = v_G2_6126_out0;
assign v_S_4421_out0 = v_G1_3852_out0;
assign v_S_4423_out0 = v_G1_3854_out0;
assign v_S_4427_out0 = v_G1_3858_out0;
assign v_S_4429_out0 = v_G1_3860_out0;
assign v_S_4431_out0 = v_G1_3862_out0;
assign v_S_4434_out0 = v_G1_3865_out0;
assign v_S_4436_out0 = v_G1_3867_out0;
assign v_S_4438_out0 = v_G1_3869_out0;
assign v_S_4440_out0 = v_G1_3871_out0;
assign v_S_4442_out0 = v_G1_3873_out0;
assign v_S_4444_out0 = v_G1_3875_out0;
assign v_S_4446_out0 = v_G1_3877_out0;
assign v_S_4448_out0 = v_G1_3879_out0;
assign v_S_4450_out0 = v_G1_3881_out0;
assign v_CIN_4870_out0 = v_CARRY_2446_out0;
assign v_MUX1_5302_out0 = v_G14_578_out0 ? v_JUMPADRESS_2316_out0 : v_REG1_210_out0;
assign v__841_out0 = { v__1570_out0,v_S_2280_out0 };
assign v_RD_2951_out0 = v_CIN_4870_out0;
assign {v_A1_3446_out1,v_A1_3446_out0 } = v_MUX1_5302_out0 + v_ADDER_IN_5411_out0 + v_G11_6620_out0;
assign v_RM_5625_out0 = v_S_4421_out0;
assign v_RM_5627_out0 = v_S_4423_out0;
assign v_RM_5631_out0 = v_S_4427_out0;
assign v_RM_5633_out0 = v_S_4429_out0;
assign v_RM_5635_out0 = v_S_4431_out0;
assign v_RM_5638_out0 = v_S_4434_out0;
assign v_RM_5640_out0 = v_S_4436_out0;
assign v_RM_5642_out0 = v_S_4438_out0;
assign v_RM_5644_out0 = v_S_4440_out0;
assign v_RM_5646_out0 = v_S_4442_out0;
assign v_RM_5648_out0 = v_S_4444_out0;
assign v_RM_5650_out0 = v_S_4446_out0;
assign v_RM_5652_out0 = v_S_4448_out0;
assign v_RM_5654_out0 = v_S_4450_out0;
assign v_COUT_36_out0 = v_A1_3446_out1;
assign v_MUX4_1295_out0 = v_BYTE_READY_1393_out0 ? v_C1_1182_out0 : v_A1_3446_out0;
assign v_G1_3870_out0 = ((v_RD_2951_out0 && !v_RM_5642_out0) || (!v_RD_2951_out0) && v_RM_5642_out0);
assign v_MUX3_5092_out0 = v_STP_5531_out0 ? v_A1_3446_out0 : v_MUX1_5302_out0;
assign v_G2_6115_out0 = v_RD_2951_out0 && v_RM_5642_out0;
assign v_CARRY_2452_out0 = v_G2_6115_out0;
assign v_PC_COUNTER_NEXT_3468_out0 = v_MUX3_5092_out0;
assign v_S_4439_out0 = v_G1_3870_out0;
assign v_PC_COUNTER_16_out0 = v_PC_COUNTER_NEXT_3468_out0;
assign v_S_634_out0 = v_S_4439_out0;
assign v_MUX1_1169_out0 = v_EXEC1LS_3338_out0 ? v_RAMADDRESSMUX_3375_out0 : v_PC_COUNTER_NEXT_3468_out0;
assign v_G1_1986_out0 = v_CARRY_2452_out0 || v_CARRY_2451_out0;
assign v_COUT_370_out0 = v_G1_1986_out0;
assign v_MUX3_1571_out0 = v_BYTE_READY_3447_out0 ? v_C2_5297_out0 : v_MUX1_1169_out0;
assign v__4281_out0 = { v_PC_COUNTER_16_out0,v_C1_980_out0 };
assign v_MUX2_1561_out0 = v_BYTE_READY_3447_out0 ? v__4281_out0 : v_RAM_IN_116_out0;
assign v_CIN_4876_out0 = v_COUT_370_out0;
assign v_NEXTADD_5180_out0 = v_MUX3_1571_out0;
assign v_NEXTADRESS_882_out0 = v_NEXTADD_5180_out0;
assign v_RD_2963_out0 = v_CIN_4876_out0;
assign v_G1_3882_out0 = ((v_RD_2963_out0 && !v_RM_5654_out0) || (!v_RD_2963_out0) && v_RM_5654_out0);
assign v_G2_6127_out0 = v_RD_2963_out0 && v_RM_5654_out0;
assign v_CARRY_2464_out0 = v_G2_6127_out0;
assign v_S_4451_out0 = v_G1_3882_out0;
assign v_S_640_out0 = v_S_4451_out0;
assign v_G1_1992_out0 = v_CARRY_2464_out0 || v_CARRY_2463_out0;
assign v_COUT_376_out0 = v_G1_1992_out0;
assign v__2337_out0 = { v_S_634_out0,v_S_640_out0 };
assign v_CIN_4871_out0 = v_COUT_376_out0;
assign v_RD_2953_out0 = v_CIN_4871_out0;
assign v_G1_3872_out0 = ((v_RD_2953_out0 && !v_RM_5644_out0) || (!v_RD_2953_out0) && v_RM_5644_out0);
assign v_G2_6117_out0 = v_RD_2953_out0 && v_RM_5644_out0;
assign v_CARRY_2454_out0 = v_G2_6117_out0;
assign v_S_4441_out0 = v_G1_3872_out0;
assign v_S_635_out0 = v_S_4441_out0;
assign v_G1_1987_out0 = v_CARRY_2454_out0 || v_CARRY_2453_out0;
assign v_COUT_371_out0 = v_G1_1987_out0;
assign v__1246_out0 = { v__2337_out0,v_S_635_out0 };
assign v_CIN_4866_out0 = v_COUT_371_out0;
assign v_RD_2942_out0 = v_CIN_4866_out0;
assign v_G1_3861_out0 = ((v_RD_2942_out0 && !v_RM_5633_out0) || (!v_RD_2942_out0) && v_RM_5633_out0);
assign v_G2_6106_out0 = v_RD_2942_out0 && v_RM_5633_out0;
assign v_CARRY_2443_out0 = v_G2_6106_out0;
assign v_S_4430_out0 = v_G1_3861_out0;
assign v_S_630_out0 = v_S_4430_out0;
assign v_G1_1982_out0 = v_CARRY_2443_out0 || v_CARRY_2442_out0;
assign v_COUT_366_out0 = v_G1_1982_out0;
assign v__3454_out0 = { v__1246_out0,v_S_630_out0 };
assign v_CIN_4865_out0 = v_COUT_366_out0;
assign v_RD_2940_out0 = v_CIN_4865_out0;
assign v_G1_3859_out0 = ((v_RD_2940_out0 && !v_RM_5631_out0) || (!v_RD_2940_out0) && v_RM_5631_out0);
assign v_G2_6104_out0 = v_RD_2940_out0 && v_RM_5631_out0;
assign v_CARRY_2441_out0 = v_G2_6104_out0;
assign v_S_4428_out0 = v_G1_3859_out0;
assign v_S_629_out0 = v_S_4428_out0;
assign v_G1_1981_out0 = v_CARRY_2441_out0 || v_CARRY_2440_out0;
assign v_COUT_365_out0 = v_G1_1981_out0;
assign v__6664_out0 = { v__3454_out0,v_S_629_out0 };
assign v_CIN_4872_out0 = v_COUT_365_out0;
assign v_RD_2955_out0 = v_CIN_4872_out0;
assign v_G1_3874_out0 = ((v_RD_2955_out0 && !v_RM_5646_out0) || (!v_RD_2955_out0) && v_RM_5646_out0);
assign v_G2_6119_out0 = v_RD_2955_out0 && v_RM_5646_out0;
assign v_CARRY_2456_out0 = v_G2_6119_out0;
assign v_S_4443_out0 = v_G1_3874_out0;
assign v_S_636_out0 = v_S_4443_out0;
assign v_G1_1988_out0 = v_CARRY_2456_out0 || v_CARRY_2455_out0;
assign v_COUT_372_out0 = v_G1_1988_out0;
assign v__1612_out0 = { v__6664_out0,v_S_636_out0 };
assign v_CIN_4873_out0 = v_COUT_372_out0;
assign v_RD_2957_out0 = v_CIN_4873_out0;
assign v_G1_3876_out0 = ((v_RD_2957_out0 && !v_RM_5648_out0) || (!v_RD_2957_out0) && v_RM_5648_out0);
assign v_G2_6121_out0 = v_RD_2957_out0 && v_RM_5648_out0;
assign v_CARRY_2458_out0 = v_G2_6121_out0;
assign v_S_4445_out0 = v_G1_3876_out0;
assign v_S_637_out0 = v_S_4445_out0;
assign v_G1_1989_out0 = v_CARRY_2458_out0 || v_CARRY_2457_out0;
assign v_COUT_373_out0 = v_G1_1989_out0;
assign v__3509_out0 = { v__1612_out0,v_S_637_out0 };
assign v_CIN_4875_out0 = v_COUT_373_out0;
assign v_RD_2961_out0 = v_CIN_4875_out0;
assign v_G1_3880_out0 = ((v_RD_2961_out0 && !v_RM_5652_out0) || (!v_RD_2961_out0) && v_RM_5652_out0);
assign v_G2_6125_out0 = v_RD_2961_out0 && v_RM_5652_out0;
assign v_CARRY_2462_out0 = v_G2_6125_out0;
assign v_S_4449_out0 = v_G1_3880_out0;
assign v_S_639_out0 = v_S_4449_out0;
assign v_G1_1991_out0 = v_CARRY_2462_out0 || v_CARRY_2461_out0;
assign v_COUT_375_out0 = v_G1_1991_out0;
assign v__2320_out0 = { v__3509_out0,v_S_639_out0 };
assign v_CIN_4868_out0 = v_COUT_375_out0;
assign v_RD_2947_out0 = v_CIN_4868_out0;
assign v_G1_3866_out0 = ((v_RD_2947_out0 && !v_RM_5638_out0) || (!v_RD_2947_out0) && v_RM_5638_out0);
assign v_G2_6111_out0 = v_RD_2947_out0 && v_RM_5638_out0;
assign v_CARRY_2448_out0 = v_G2_6111_out0;
assign v_S_4435_out0 = v_G1_3866_out0;
assign v_S_632_out0 = v_S_4435_out0;
assign v_G1_1984_out0 = v_CARRY_2448_out0 || v_CARRY_2447_out0;
assign v_COUT_368_out0 = v_G1_1984_out0;
assign v__3402_out0 = { v__2320_out0,v_S_632_out0 };
assign v_CIN_4869_out0 = v_COUT_368_out0;
assign v_RD_2949_out0 = v_CIN_4869_out0;
assign v_G1_3868_out0 = ((v_RD_2949_out0 && !v_RM_5640_out0) || (!v_RD_2949_out0) && v_RM_5640_out0);
assign v_G2_6113_out0 = v_RD_2949_out0 && v_RM_5640_out0;
assign v_CARRY_2450_out0 = v_G2_6113_out0;
assign v_S_4437_out0 = v_G1_3868_out0;
assign v_S_633_out0 = v_S_4437_out0;
assign v_G1_1985_out0 = v_CARRY_2450_out0 || v_CARRY_2449_out0;
assign v_COUT_369_out0 = v_G1_1985_out0;
assign v__2846_out0 = { v__3402_out0,v_S_633_out0 };
assign v_CIN_4874_out0 = v_COUT_369_out0;
assign v_RD_2959_out0 = v_CIN_4874_out0;
assign v_G1_3878_out0 = ((v_RD_2959_out0 && !v_RM_5650_out0) || (!v_RD_2959_out0) && v_RM_5650_out0);
assign v_G2_6123_out0 = v_RD_2959_out0 && v_RM_5650_out0;
assign v_CARRY_2460_out0 = v_G2_6123_out0;
assign v_S_4447_out0 = v_G1_3878_out0;
assign v_S_638_out0 = v_S_4447_out0;
assign v_G1_1990_out0 = v_CARRY_2460_out0 || v_CARRY_2459_out0;
assign v_COUT_374_out0 = v_G1_1990_out0;
assign v__990_out0 = { v__2846_out0,v_S_638_out0 };
assign v_CIN_4862_out0 = v_COUT_374_out0;
assign v_RD_2934_out0 = v_CIN_4862_out0;
assign v_G1_3853_out0 = ((v_RD_2934_out0 && !v_RM_5625_out0) || (!v_RD_2934_out0) && v_RM_5625_out0);
assign v_G2_6098_out0 = v_RD_2934_out0 && v_RM_5625_out0;
assign v_CARRY_2435_out0 = v_G2_6098_out0;
assign v_S_4422_out0 = v_G1_3853_out0;
assign v_S_626_out0 = v_S_4422_out0;
assign v_G1_1978_out0 = v_CARRY_2435_out0 || v_CARRY_2434_out0;
assign v_COUT_362_out0 = v_G1_1978_out0;
assign v__1366_out0 = { v__990_out0,v_S_626_out0 };
assign v_CIN_4867_out0 = v_COUT_362_out0;
assign v_RD_2944_out0 = v_CIN_4867_out0;
assign v_G1_3863_out0 = ((v_RD_2944_out0 && !v_RM_5635_out0) || (!v_RD_2944_out0) && v_RM_5635_out0);
assign v_G2_6108_out0 = v_RD_2944_out0 && v_RM_5635_out0;
assign v_CARRY_2445_out0 = v_G2_6108_out0;
assign v_S_4432_out0 = v_G1_3863_out0;
assign v_S_631_out0 = v_S_4432_out0;
assign v_G1_1983_out0 = v_CARRY_2445_out0 || v_CARRY_2444_out0;
assign v_COUT_367_out0 = v_G1_1983_out0;
assign v__893_out0 = { v__1366_out0,v_S_631_out0 };
assign v_CIN_4863_out0 = v_COUT_367_out0;
assign v_RD_2936_out0 = v_CIN_4863_out0;
assign v_G1_3855_out0 = ((v_RD_2936_out0 && !v_RM_5627_out0) || (!v_RD_2936_out0) && v_RM_5627_out0);
assign v_G2_6100_out0 = v_RD_2936_out0 && v_RM_5627_out0;
assign v_CARRY_2437_out0 = v_G2_6100_out0;
assign v_S_4424_out0 = v_G1_3855_out0;
assign v_S_627_out0 = v_S_4424_out0;
assign v_G1_1979_out0 = v_CARRY_2437_out0 || v_CARRY_2436_out0;
assign v_COUT_363_out0 = v_G1_1979_out0;
assign v__2222_out0 = { v__893_out0,v_S_627_out0 };
assign v_RM_1661_out0 = v_COUT_363_out0;
assign v_RM_5628_out0 = v_RM_1661_out0;
assign v_G1_3856_out0 = ((v_RD_2937_out0 && !v_RM_5628_out0) || (!v_RD_2937_out0) && v_RM_5628_out0);
assign v_G2_6101_out0 = v_RD_2937_out0 && v_RM_5628_out0;
assign v_CARRY_2438_out0 = v_G2_6101_out0;
assign v_S_4425_out0 = v_G1_3856_out0;
assign v_RM_5629_out0 = v_S_4425_out0;
assign v_G1_3857_out0 = ((v_RD_2938_out0 && !v_RM_5629_out0) || (!v_RD_2938_out0) && v_RM_5629_out0);
assign v_G2_6102_out0 = v_RD_2938_out0 && v_RM_5629_out0;
assign v_CARRY_2439_out0 = v_G2_6102_out0;
assign v_S_4426_out0 = v_G1_3857_out0;
assign v_S_628_out0 = v_S_4426_out0;
assign v_G1_1980_out0 = v_CARRY_2439_out0 || v_CARRY_2438_out0;
assign v_COUT_364_out0 = v_G1_1980_out0;
assign v__5245_out0 = { v__2222_out0,v_S_628_out0 };
assign v__5388_out0 = { v__5245_out0,v_COUT_364_out0 };
assign v_COUT_5373_out0 = v__5388_out0;
assign v_CIN_1151_out0 = v_COUT_5373_out0;
assign v__233_out0 = v_CIN_1151_out0[8:8];
assign v__871_out0 = v_CIN_1151_out0[6:6];
assign v__1054_out0 = v_CIN_1151_out0[3:3];
assign v__1073_out0 = v_CIN_1151_out0[15:15];
assign v__1224_out0 = v_CIN_1151_out0[0:0];
assign v__1492_out0 = v_CIN_1151_out0[9:9];
assign v__1508_out0 = v_CIN_1151_out0[2:2];
assign v__1534_out0 = v_CIN_1151_out0[7:7];
assign v__1867_out0 = v_CIN_1151_out0[1:1];
assign v__1885_out0 = v_CIN_1151_out0[10:10];
assign v__3344_out0 = v_CIN_1151_out0[11:11];
assign v__3760_out0 = v_CIN_1151_out0[12:12];
assign v__4286_out0 = v_CIN_1151_out0[13:13];
assign v__4319_out0 = v_CIN_1151_out0[14:14];
assign v__5280_out0 = v_CIN_1151_out0[5:5];
assign v__6628_out0 = v_CIN_1151_out0[4:4];
assign v_RM_1689_out0 = v__3760_out0;
assign v_RM_1690_out0 = v__4319_out0;
assign v_RM_1692_out0 = v__5280_out0;
assign v_RM_1693_out0 = v__6628_out0;
assign v_RM_1694_out0 = v__4286_out0;
assign v_RM_1695_out0 = v__1492_out0;
assign v_RM_1696_out0 = v__1885_out0;
assign v_RM_1697_out0 = v__1867_out0;
assign v_RM_1698_out0 = v__1054_out0;
assign v_RM_1699_out0 = v__871_out0;
assign v_RM_1700_out0 = v__1534_out0;
assign v_RM_1701_out0 = v__3344_out0;
assign v_RM_1702_out0 = v__233_out0;
assign v_RM_1703_out0 = v__1508_out0;
assign v_CIN_4894_out0 = v__1073_out0;
assign v_RM_5698_out0 = v__1224_out0;
assign v_RD_3000_out0 = v_CIN_4894_out0;
assign v_G1_3926_out0 = ((v_RD_3007_out0 && !v_RM_5698_out0) || (!v_RD_3007_out0) && v_RM_5698_out0);
assign v_RM_5686_out0 = v_RM_1689_out0;
assign v_RM_5688_out0 = v_RM_1690_out0;
assign v_RM_5692_out0 = v_RM_1692_out0;
assign v_RM_5694_out0 = v_RM_1693_out0;
assign v_RM_5696_out0 = v_RM_1694_out0;
assign v_RM_5699_out0 = v_RM_1695_out0;
assign v_RM_5701_out0 = v_RM_1696_out0;
assign v_RM_5703_out0 = v_RM_1697_out0;
assign v_RM_5705_out0 = v_RM_1698_out0;
assign v_RM_5707_out0 = v_RM_1699_out0;
assign v_RM_5709_out0 = v_RM_1700_out0;
assign v_RM_5711_out0 = v_RM_1701_out0;
assign v_RM_5713_out0 = v_RM_1702_out0;
assign v_RM_5715_out0 = v_RM_1703_out0;
assign v_G2_6171_out0 = v_RD_3007_out0 && v_RM_5698_out0;
assign v_CARRY_2508_out0 = v_G2_6171_out0;
assign v_G1_3914_out0 = ((v_RD_2995_out0 && !v_RM_5686_out0) || (!v_RD_2995_out0) && v_RM_5686_out0);
assign v_G1_3916_out0 = ((v_RD_2997_out0 && !v_RM_5688_out0) || (!v_RD_2997_out0) && v_RM_5688_out0);
assign v_G1_3920_out0 = ((v_RD_3001_out0 && !v_RM_5692_out0) || (!v_RD_3001_out0) && v_RM_5692_out0);
assign v_G1_3922_out0 = ((v_RD_3003_out0 && !v_RM_5694_out0) || (!v_RD_3003_out0) && v_RM_5694_out0);
assign v_G1_3924_out0 = ((v_RD_3005_out0 && !v_RM_5696_out0) || (!v_RD_3005_out0) && v_RM_5696_out0);
assign v_G1_3927_out0 = ((v_RD_3008_out0 && !v_RM_5699_out0) || (!v_RD_3008_out0) && v_RM_5699_out0);
assign v_G1_3929_out0 = ((v_RD_3010_out0 && !v_RM_5701_out0) || (!v_RD_3010_out0) && v_RM_5701_out0);
assign v_G1_3931_out0 = ((v_RD_3012_out0 && !v_RM_5703_out0) || (!v_RD_3012_out0) && v_RM_5703_out0);
assign v_G1_3933_out0 = ((v_RD_3014_out0 && !v_RM_5705_out0) || (!v_RD_3014_out0) && v_RM_5705_out0);
assign v_G1_3935_out0 = ((v_RD_3016_out0 && !v_RM_5707_out0) || (!v_RD_3016_out0) && v_RM_5707_out0);
assign v_G1_3937_out0 = ((v_RD_3018_out0 && !v_RM_5709_out0) || (!v_RD_3018_out0) && v_RM_5709_out0);
assign v_G1_3939_out0 = ((v_RD_3020_out0 && !v_RM_5711_out0) || (!v_RD_3020_out0) && v_RM_5711_out0);
assign v_G1_3941_out0 = ((v_RD_3022_out0 && !v_RM_5713_out0) || (!v_RD_3022_out0) && v_RM_5713_out0);
assign v_G1_3943_out0 = ((v_RD_3024_out0 && !v_RM_5715_out0) || (!v_RD_3024_out0) && v_RM_5715_out0);
assign v_S_4495_out0 = v_G1_3926_out0;
assign v_G2_6159_out0 = v_RD_2995_out0 && v_RM_5686_out0;
assign v_G2_6161_out0 = v_RD_2997_out0 && v_RM_5688_out0;
assign v_G2_6165_out0 = v_RD_3001_out0 && v_RM_5692_out0;
assign v_G2_6167_out0 = v_RD_3003_out0 && v_RM_5694_out0;
assign v_G2_6169_out0 = v_RD_3005_out0 && v_RM_5696_out0;
assign v_G2_6172_out0 = v_RD_3008_out0 && v_RM_5699_out0;
assign v_G2_6174_out0 = v_RD_3010_out0 && v_RM_5701_out0;
assign v_G2_6176_out0 = v_RD_3012_out0 && v_RM_5703_out0;
assign v_G2_6178_out0 = v_RD_3014_out0 && v_RM_5705_out0;
assign v_G2_6180_out0 = v_RD_3016_out0 && v_RM_5707_out0;
assign v_G2_6182_out0 = v_RD_3018_out0 && v_RM_5709_out0;
assign v_G2_6184_out0 = v_RD_3020_out0 && v_RM_5711_out0;
assign v_G2_6186_out0 = v_RD_3022_out0 && v_RM_5713_out0;
assign v_G2_6188_out0 = v_RD_3024_out0 && v_RM_5715_out0;
assign v_S_2282_out0 = v_S_4495_out0;
assign v_CARRY_2496_out0 = v_G2_6159_out0;
assign v_CARRY_2498_out0 = v_G2_6161_out0;
assign v_CARRY_2502_out0 = v_G2_6165_out0;
assign v_CARRY_2504_out0 = v_G2_6167_out0;
assign v_CARRY_2506_out0 = v_G2_6169_out0;
assign v_CARRY_2509_out0 = v_G2_6172_out0;
assign v_CARRY_2511_out0 = v_G2_6174_out0;
assign v_CARRY_2513_out0 = v_G2_6176_out0;
assign v_CARRY_2515_out0 = v_G2_6178_out0;
assign v_CARRY_2517_out0 = v_G2_6180_out0;
assign v_CARRY_2519_out0 = v_G2_6182_out0;
assign v_CARRY_2521_out0 = v_G2_6184_out0;
assign v_CARRY_2523_out0 = v_G2_6186_out0;
assign v_CARRY_2525_out0 = v_G2_6188_out0;
assign v_S_4483_out0 = v_G1_3914_out0;
assign v_S_4485_out0 = v_G1_3916_out0;
assign v_S_4489_out0 = v_G1_3920_out0;
assign v_S_4491_out0 = v_G1_3922_out0;
assign v_S_4493_out0 = v_G1_3924_out0;
assign v_S_4496_out0 = v_G1_3927_out0;
assign v_S_4498_out0 = v_G1_3929_out0;
assign v_S_4500_out0 = v_G1_3931_out0;
assign v_S_4502_out0 = v_G1_3933_out0;
assign v_S_4504_out0 = v_G1_3935_out0;
assign v_S_4506_out0 = v_G1_3937_out0;
assign v_S_4508_out0 = v_G1_3939_out0;
assign v_S_4510_out0 = v_G1_3941_out0;
assign v_S_4512_out0 = v_G1_3943_out0;
assign v_CIN_4900_out0 = v_CARRY_2508_out0;
assign v__2213_out0 = { v__841_out0,v_S_2282_out0 };
assign v_RD_3013_out0 = v_CIN_4900_out0;
assign v_RM_5687_out0 = v_S_4483_out0;
assign v_RM_5689_out0 = v_S_4485_out0;
assign v_RM_5693_out0 = v_S_4489_out0;
assign v_RM_5695_out0 = v_S_4491_out0;
assign v_RM_5697_out0 = v_S_4493_out0;
assign v_RM_5700_out0 = v_S_4496_out0;
assign v_RM_5702_out0 = v_S_4498_out0;
assign v_RM_5704_out0 = v_S_4500_out0;
assign v_RM_5706_out0 = v_S_4502_out0;
assign v_RM_5708_out0 = v_S_4504_out0;
assign v_RM_5710_out0 = v_S_4506_out0;
assign v_RM_5712_out0 = v_S_4508_out0;
assign v_RM_5714_out0 = v_S_4510_out0;
assign v_RM_5716_out0 = v_S_4512_out0;
assign v_G1_3932_out0 = ((v_RD_3013_out0 && !v_RM_5704_out0) || (!v_RD_3013_out0) && v_RM_5704_out0);
assign v_G2_6177_out0 = v_RD_3013_out0 && v_RM_5704_out0;
assign v_CARRY_2514_out0 = v_G2_6177_out0;
assign v_S_4501_out0 = v_G1_3932_out0;
assign v_S_664_out0 = v_S_4501_out0;
assign v_G1_2016_out0 = v_CARRY_2514_out0 || v_CARRY_2513_out0;
assign v_COUT_400_out0 = v_G1_2016_out0;
assign v_CIN_4906_out0 = v_COUT_400_out0;
assign v_RD_3025_out0 = v_CIN_4906_out0;
assign v_G1_3944_out0 = ((v_RD_3025_out0 && !v_RM_5716_out0) || (!v_RD_3025_out0) && v_RM_5716_out0);
assign v_G2_6189_out0 = v_RD_3025_out0 && v_RM_5716_out0;
assign v_CARRY_2526_out0 = v_G2_6189_out0;
assign v_S_4513_out0 = v_G1_3944_out0;
assign v_S_670_out0 = v_S_4513_out0;
assign v_G1_2022_out0 = v_CARRY_2526_out0 || v_CARRY_2525_out0;
assign v_COUT_406_out0 = v_G1_2022_out0;
assign v__2339_out0 = { v_S_664_out0,v_S_670_out0 };
assign v_CIN_4901_out0 = v_COUT_406_out0;
assign v_RD_3015_out0 = v_CIN_4901_out0;
assign v_G1_3934_out0 = ((v_RD_3015_out0 && !v_RM_5706_out0) || (!v_RD_3015_out0) && v_RM_5706_out0);
assign v_G2_6179_out0 = v_RD_3015_out0 && v_RM_5706_out0;
assign v_CARRY_2516_out0 = v_G2_6179_out0;
assign v_S_4503_out0 = v_G1_3934_out0;
assign v_S_665_out0 = v_S_4503_out0;
assign v_G1_2017_out0 = v_CARRY_2516_out0 || v_CARRY_2515_out0;
assign v_COUT_401_out0 = v_G1_2017_out0;
assign v__1248_out0 = { v__2339_out0,v_S_665_out0 };
assign v_CIN_4896_out0 = v_COUT_401_out0;
assign v_RD_3004_out0 = v_CIN_4896_out0;
assign v_G1_3923_out0 = ((v_RD_3004_out0 && !v_RM_5695_out0) || (!v_RD_3004_out0) && v_RM_5695_out0);
assign v_G2_6168_out0 = v_RD_3004_out0 && v_RM_5695_out0;
assign v_CARRY_2505_out0 = v_G2_6168_out0;
assign v_S_4492_out0 = v_G1_3923_out0;
assign v_S_660_out0 = v_S_4492_out0;
assign v_G1_2012_out0 = v_CARRY_2505_out0 || v_CARRY_2504_out0;
assign v_COUT_396_out0 = v_G1_2012_out0;
assign v__3456_out0 = { v__1248_out0,v_S_660_out0 };
assign v_CIN_4895_out0 = v_COUT_396_out0;
assign v_RD_3002_out0 = v_CIN_4895_out0;
assign v_G1_3921_out0 = ((v_RD_3002_out0 && !v_RM_5693_out0) || (!v_RD_3002_out0) && v_RM_5693_out0);
assign v_G2_6166_out0 = v_RD_3002_out0 && v_RM_5693_out0;
assign v_CARRY_2503_out0 = v_G2_6166_out0;
assign v_S_4490_out0 = v_G1_3921_out0;
assign v_S_659_out0 = v_S_4490_out0;
assign v_G1_2011_out0 = v_CARRY_2503_out0 || v_CARRY_2502_out0;
assign v_COUT_395_out0 = v_G1_2011_out0;
assign v__6666_out0 = { v__3456_out0,v_S_659_out0 };
assign v_CIN_4902_out0 = v_COUT_395_out0;
assign v_RD_3017_out0 = v_CIN_4902_out0;
assign v_G1_3936_out0 = ((v_RD_3017_out0 && !v_RM_5708_out0) || (!v_RD_3017_out0) && v_RM_5708_out0);
assign v_G2_6181_out0 = v_RD_3017_out0 && v_RM_5708_out0;
assign v_CARRY_2518_out0 = v_G2_6181_out0;
assign v_S_4505_out0 = v_G1_3936_out0;
assign v_S_666_out0 = v_S_4505_out0;
assign v_G1_2018_out0 = v_CARRY_2518_out0 || v_CARRY_2517_out0;
assign v_COUT_402_out0 = v_G1_2018_out0;
assign v__1614_out0 = { v__6666_out0,v_S_666_out0 };
assign v_CIN_4903_out0 = v_COUT_402_out0;
assign v_RD_3019_out0 = v_CIN_4903_out0;
assign v_G1_3938_out0 = ((v_RD_3019_out0 && !v_RM_5710_out0) || (!v_RD_3019_out0) && v_RM_5710_out0);
assign v_G2_6183_out0 = v_RD_3019_out0 && v_RM_5710_out0;
assign v_CARRY_2520_out0 = v_G2_6183_out0;
assign v_S_4507_out0 = v_G1_3938_out0;
assign v_S_667_out0 = v_S_4507_out0;
assign v_G1_2019_out0 = v_CARRY_2520_out0 || v_CARRY_2519_out0;
assign v_COUT_403_out0 = v_G1_2019_out0;
assign v__3511_out0 = { v__1614_out0,v_S_667_out0 };
assign v_CIN_4905_out0 = v_COUT_403_out0;
assign v_RD_3023_out0 = v_CIN_4905_out0;
assign v_G1_3942_out0 = ((v_RD_3023_out0 && !v_RM_5714_out0) || (!v_RD_3023_out0) && v_RM_5714_out0);
assign v_G2_6187_out0 = v_RD_3023_out0 && v_RM_5714_out0;
assign v_CARRY_2524_out0 = v_G2_6187_out0;
assign v_S_4511_out0 = v_G1_3942_out0;
assign v_S_669_out0 = v_S_4511_out0;
assign v_G1_2021_out0 = v_CARRY_2524_out0 || v_CARRY_2523_out0;
assign v_COUT_405_out0 = v_G1_2021_out0;
assign v__2322_out0 = { v__3511_out0,v_S_669_out0 };
assign v_CIN_4898_out0 = v_COUT_405_out0;
assign v_RD_3009_out0 = v_CIN_4898_out0;
assign v_G1_3928_out0 = ((v_RD_3009_out0 && !v_RM_5700_out0) || (!v_RD_3009_out0) && v_RM_5700_out0);
assign v_G2_6173_out0 = v_RD_3009_out0 && v_RM_5700_out0;
assign v_CARRY_2510_out0 = v_G2_6173_out0;
assign v_S_4497_out0 = v_G1_3928_out0;
assign v_S_662_out0 = v_S_4497_out0;
assign v_G1_2014_out0 = v_CARRY_2510_out0 || v_CARRY_2509_out0;
assign v_COUT_398_out0 = v_G1_2014_out0;
assign v__3404_out0 = { v__2322_out0,v_S_662_out0 };
assign v_CIN_4899_out0 = v_COUT_398_out0;
assign v_RD_3011_out0 = v_CIN_4899_out0;
assign v_G1_3930_out0 = ((v_RD_3011_out0 && !v_RM_5702_out0) || (!v_RD_3011_out0) && v_RM_5702_out0);
assign v_G2_6175_out0 = v_RD_3011_out0 && v_RM_5702_out0;
assign v_CARRY_2512_out0 = v_G2_6175_out0;
assign v_S_4499_out0 = v_G1_3930_out0;
assign v_S_663_out0 = v_S_4499_out0;
assign v_G1_2015_out0 = v_CARRY_2512_out0 || v_CARRY_2511_out0;
assign v_COUT_399_out0 = v_G1_2015_out0;
assign v__2848_out0 = { v__3404_out0,v_S_663_out0 };
assign v_CIN_4904_out0 = v_COUT_399_out0;
assign v_RD_3021_out0 = v_CIN_4904_out0;
assign v_G1_3940_out0 = ((v_RD_3021_out0 && !v_RM_5712_out0) || (!v_RD_3021_out0) && v_RM_5712_out0);
assign v_G2_6185_out0 = v_RD_3021_out0 && v_RM_5712_out0;
assign v_CARRY_2522_out0 = v_G2_6185_out0;
assign v_S_4509_out0 = v_G1_3940_out0;
assign v_S_668_out0 = v_S_4509_out0;
assign v_G1_2020_out0 = v_CARRY_2522_out0 || v_CARRY_2521_out0;
assign v_COUT_404_out0 = v_G1_2020_out0;
assign v__992_out0 = { v__2848_out0,v_S_668_out0 };
assign v_CIN_4892_out0 = v_COUT_404_out0;
assign v_RD_2996_out0 = v_CIN_4892_out0;
assign v_G1_3915_out0 = ((v_RD_2996_out0 && !v_RM_5687_out0) || (!v_RD_2996_out0) && v_RM_5687_out0);
assign v_G2_6160_out0 = v_RD_2996_out0 && v_RM_5687_out0;
assign v_CARRY_2497_out0 = v_G2_6160_out0;
assign v_S_4484_out0 = v_G1_3915_out0;
assign v_S_656_out0 = v_S_4484_out0;
assign v_G1_2008_out0 = v_CARRY_2497_out0 || v_CARRY_2496_out0;
assign v_COUT_392_out0 = v_G1_2008_out0;
assign v__1368_out0 = { v__992_out0,v_S_656_out0 };
assign v_CIN_4897_out0 = v_COUT_392_out0;
assign v_RD_3006_out0 = v_CIN_4897_out0;
assign v_G1_3925_out0 = ((v_RD_3006_out0 && !v_RM_5697_out0) || (!v_RD_3006_out0) && v_RM_5697_out0);
assign v_G2_6170_out0 = v_RD_3006_out0 && v_RM_5697_out0;
assign v_CARRY_2507_out0 = v_G2_6170_out0;
assign v_S_4494_out0 = v_G1_3925_out0;
assign v_S_661_out0 = v_S_4494_out0;
assign v_G1_2013_out0 = v_CARRY_2507_out0 || v_CARRY_2506_out0;
assign v_COUT_397_out0 = v_G1_2013_out0;
assign v__895_out0 = { v__1368_out0,v_S_661_out0 };
assign v_CIN_4893_out0 = v_COUT_397_out0;
assign v_RD_2998_out0 = v_CIN_4893_out0;
assign v_G1_3917_out0 = ((v_RD_2998_out0 && !v_RM_5689_out0) || (!v_RD_2998_out0) && v_RM_5689_out0);
assign v_G2_6162_out0 = v_RD_2998_out0 && v_RM_5689_out0;
assign v_CARRY_2499_out0 = v_G2_6162_out0;
assign v_S_4486_out0 = v_G1_3917_out0;
assign v_S_657_out0 = v_S_4486_out0;
assign v_G1_2009_out0 = v_CARRY_2499_out0 || v_CARRY_2498_out0;
assign v_COUT_393_out0 = v_G1_2009_out0;
assign v__2224_out0 = { v__895_out0,v_S_657_out0 };
assign v_RM_1691_out0 = v_COUT_393_out0;
assign v_RM_5690_out0 = v_RM_1691_out0;
assign v_G1_3918_out0 = ((v_RD_2999_out0 && !v_RM_5690_out0) || (!v_RD_2999_out0) && v_RM_5690_out0);
assign v_G2_6163_out0 = v_RD_2999_out0 && v_RM_5690_out0;
assign v_CARRY_2500_out0 = v_G2_6163_out0;
assign v_S_4487_out0 = v_G1_3918_out0;
assign v_RM_5691_out0 = v_S_4487_out0;
assign v_G1_3919_out0 = ((v_RD_3000_out0 && !v_RM_5691_out0) || (!v_RD_3000_out0) && v_RM_5691_out0);
assign v_G2_6164_out0 = v_RD_3000_out0 && v_RM_5691_out0;
assign v_CARRY_2501_out0 = v_G2_6164_out0;
assign v_S_4488_out0 = v_G1_3919_out0;
assign v_S_658_out0 = v_S_4488_out0;
assign v_G1_2010_out0 = v_CARRY_2501_out0 || v_CARRY_2500_out0;
assign v_COUT_394_out0 = v_G1_2010_out0;
assign v__5247_out0 = { v__2224_out0,v_S_658_out0 };
assign v__5390_out0 = { v__5247_out0,v_COUT_394_out0 };
assign v_COUT_5375_out0 = v__5390_out0;
assign v_CIN_1147_out0 = v_COUT_5375_out0;
assign v__229_out0 = v_CIN_1147_out0[8:8];
assign v__867_out0 = v_CIN_1147_out0[6:6];
assign v__1050_out0 = v_CIN_1147_out0[3:3];
assign v__1070_out0 = v_CIN_1147_out0[15:15];
assign v__1220_out0 = v_CIN_1147_out0[0:0];
assign v__1488_out0 = v_CIN_1147_out0[9:9];
assign v__1504_out0 = v_CIN_1147_out0[2:2];
assign v__1530_out0 = v_CIN_1147_out0[7:7];
assign v__1863_out0 = v_CIN_1147_out0[1:1];
assign v__1881_out0 = v_CIN_1147_out0[10:10];
assign v__3340_out0 = v_CIN_1147_out0[11:11];
assign v__3756_out0 = v_CIN_1147_out0[12:12];
assign v__4282_out0 = v_CIN_1147_out0[13:13];
assign v__4315_out0 = v_CIN_1147_out0[14:14];
assign v__5276_out0 = v_CIN_1147_out0[5:5];
assign v__6624_out0 = v_CIN_1147_out0[4:4];
assign v_RM_1630_out0 = v__3756_out0;
assign v_RM_1631_out0 = v__4315_out0;
assign v_RM_1633_out0 = v__5276_out0;
assign v_RM_1634_out0 = v__6624_out0;
assign v_RM_1635_out0 = v__4282_out0;
assign v_RM_1636_out0 = v__1488_out0;
assign v_RM_1637_out0 = v__1881_out0;
assign v_RM_1638_out0 = v__1863_out0;
assign v_RM_1639_out0 = v__1050_out0;
assign v_RM_1640_out0 = v__867_out0;
assign v_RM_1641_out0 = v__1530_out0;
assign v_RM_1642_out0 = v__3340_out0;
assign v_RM_1643_out0 = v__229_out0;
assign v_RM_1644_out0 = v__1504_out0;
assign v_CIN_4835_out0 = v__1070_out0;
assign v_RM_5575_out0 = v__1220_out0;
assign v_RD_2877_out0 = v_CIN_4835_out0;
assign v_G1_3803_out0 = ((v_RD_2884_out0 && !v_RM_5575_out0) || (!v_RD_2884_out0) && v_RM_5575_out0);
assign v_RM_5563_out0 = v_RM_1630_out0;
assign v_RM_5565_out0 = v_RM_1631_out0;
assign v_RM_5569_out0 = v_RM_1633_out0;
assign v_RM_5571_out0 = v_RM_1634_out0;
assign v_RM_5573_out0 = v_RM_1635_out0;
assign v_RM_5576_out0 = v_RM_1636_out0;
assign v_RM_5578_out0 = v_RM_1637_out0;
assign v_RM_5580_out0 = v_RM_1638_out0;
assign v_RM_5582_out0 = v_RM_1639_out0;
assign v_RM_5584_out0 = v_RM_1640_out0;
assign v_RM_5586_out0 = v_RM_1641_out0;
assign v_RM_5588_out0 = v_RM_1642_out0;
assign v_RM_5590_out0 = v_RM_1643_out0;
assign v_RM_5592_out0 = v_RM_1644_out0;
assign v_G2_6048_out0 = v_RD_2884_out0 && v_RM_5575_out0;
assign v_CARRY_2385_out0 = v_G2_6048_out0;
assign v_G1_3791_out0 = ((v_RD_2872_out0 && !v_RM_5563_out0) || (!v_RD_2872_out0) && v_RM_5563_out0);
assign v_G1_3793_out0 = ((v_RD_2874_out0 && !v_RM_5565_out0) || (!v_RD_2874_out0) && v_RM_5565_out0);
assign v_G1_3797_out0 = ((v_RD_2878_out0 && !v_RM_5569_out0) || (!v_RD_2878_out0) && v_RM_5569_out0);
assign v_G1_3799_out0 = ((v_RD_2880_out0 && !v_RM_5571_out0) || (!v_RD_2880_out0) && v_RM_5571_out0);
assign v_G1_3801_out0 = ((v_RD_2882_out0 && !v_RM_5573_out0) || (!v_RD_2882_out0) && v_RM_5573_out0);
assign v_G1_3804_out0 = ((v_RD_2885_out0 && !v_RM_5576_out0) || (!v_RD_2885_out0) && v_RM_5576_out0);
assign v_G1_3806_out0 = ((v_RD_2887_out0 && !v_RM_5578_out0) || (!v_RD_2887_out0) && v_RM_5578_out0);
assign v_G1_3808_out0 = ((v_RD_2889_out0 && !v_RM_5580_out0) || (!v_RD_2889_out0) && v_RM_5580_out0);
assign v_G1_3810_out0 = ((v_RD_2891_out0 && !v_RM_5582_out0) || (!v_RD_2891_out0) && v_RM_5582_out0);
assign v_G1_3812_out0 = ((v_RD_2893_out0 && !v_RM_5584_out0) || (!v_RD_2893_out0) && v_RM_5584_out0);
assign v_G1_3814_out0 = ((v_RD_2895_out0 && !v_RM_5586_out0) || (!v_RD_2895_out0) && v_RM_5586_out0);
assign v_G1_3816_out0 = ((v_RD_2897_out0 && !v_RM_5588_out0) || (!v_RD_2897_out0) && v_RM_5588_out0);
assign v_G1_3818_out0 = ((v_RD_2899_out0 && !v_RM_5590_out0) || (!v_RD_2899_out0) && v_RM_5590_out0);
assign v_G1_3820_out0 = ((v_RD_2901_out0 && !v_RM_5592_out0) || (!v_RD_2901_out0) && v_RM_5592_out0);
assign v_S_4372_out0 = v_G1_3803_out0;
assign v_G2_6036_out0 = v_RD_2872_out0 && v_RM_5563_out0;
assign v_G2_6038_out0 = v_RD_2874_out0 && v_RM_5565_out0;
assign v_G2_6042_out0 = v_RD_2878_out0 && v_RM_5569_out0;
assign v_G2_6044_out0 = v_RD_2880_out0 && v_RM_5571_out0;
assign v_G2_6046_out0 = v_RD_2882_out0 && v_RM_5573_out0;
assign v_G2_6049_out0 = v_RD_2885_out0 && v_RM_5576_out0;
assign v_G2_6051_out0 = v_RD_2887_out0 && v_RM_5578_out0;
assign v_G2_6053_out0 = v_RD_2889_out0 && v_RM_5580_out0;
assign v_G2_6055_out0 = v_RD_2891_out0 && v_RM_5582_out0;
assign v_G2_6057_out0 = v_RD_2893_out0 && v_RM_5584_out0;
assign v_G2_6059_out0 = v_RD_2895_out0 && v_RM_5586_out0;
assign v_G2_6061_out0 = v_RD_2897_out0 && v_RM_5588_out0;
assign v_G2_6063_out0 = v_RD_2899_out0 && v_RM_5590_out0;
assign v_G2_6065_out0 = v_RD_2901_out0 && v_RM_5592_out0;
assign v_S_2278_out0 = v_S_4372_out0;
assign v_CARRY_2373_out0 = v_G2_6036_out0;
assign v_CARRY_2375_out0 = v_G2_6038_out0;
assign v_CARRY_2379_out0 = v_G2_6042_out0;
assign v_CARRY_2381_out0 = v_G2_6044_out0;
assign v_CARRY_2383_out0 = v_G2_6046_out0;
assign v_CARRY_2386_out0 = v_G2_6049_out0;
assign v_CARRY_2388_out0 = v_G2_6051_out0;
assign v_CARRY_2390_out0 = v_G2_6053_out0;
assign v_CARRY_2392_out0 = v_G2_6055_out0;
assign v_CARRY_2394_out0 = v_G2_6057_out0;
assign v_CARRY_2396_out0 = v_G2_6059_out0;
assign v_CARRY_2398_out0 = v_G2_6061_out0;
assign v_CARRY_2400_out0 = v_G2_6063_out0;
assign v_CARRY_2402_out0 = v_G2_6065_out0;
assign v_S_4360_out0 = v_G1_3791_out0;
assign v_S_4362_out0 = v_G1_3793_out0;
assign v_S_4366_out0 = v_G1_3797_out0;
assign v_S_4368_out0 = v_G1_3799_out0;
assign v_S_4370_out0 = v_G1_3801_out0;
assign v_S_4373_out0 = v_G1_3804_out0;
assign v_S_4375_out0 = v_G1_3806_out0;
assign v_S_4377_out0 = v_G1_3808_out0;
assign v_S_4379_out0 = v_G1_3810_out0;
assign v_S_4381_out0 = v_G1_3812_out0;
assign v_S_4383_out0 = v_G1_3814_out0;
assign v_S_4385_out0 = v_G1_3816_out0;
assign v_S_4387_out0 = v_G1_3818_out0;
assign v_S_4389_out0 = v_G1_3820_out0;
assign v_CIN_4841_out0 = v_CARRY_2385_out0;
assign v__1166_out0 = { v__2213_out0,v_S_2278_out0 };
assign v_RD_2890_out0 = v_CIN_4841_out0;
assign v_RM_5564_out0 = v_S_4360_out0;
assign v_RM_5566_out0 = v_S_4362_out0;
assign v_RM_5570_out0 = v_S_4366_out0;
assign v_RM_5572_out0 = v_S_4368_out0;
assign v_RM_5574_out0 = v_S_4370_out0;
assign v_RM_5577_out0 = v_S_4373_out0;
assign v_RM_5579_out0 = v_S_4375_out0;
assign v_RM_5581_out0 = v_S_4377_out0;
assign v_RM_5583_out0 = v_S_4379_out0;
assign v_RM_5585_out0 = v_S_4381_out0;
assign v_RM_5587_out0 = v_S_4383_out0;
assign v_RM_5589_out0 = v_S_4385_out0;
assign v_RM_5591_out0 = v_S_4387_out0;
assign v_RM_5593_out0 = v_S_4389_out0;
assign v_G1_3809_out0 = ((v_RD_2890_out0 && !v_RM_5581_out0) || (!v_RD_2890_out0) && v_RM_5581_out0);
assign v_G2_6054_out0 = v_RD_2890_out0 && v_RM_5581_out0;
assign v_CARRY_2391_out0 = v_G2_6054_out0;
assign v_S_4378_out0 = v_G1_3809_out0;
assign v_S_605_out0 = v_S_4378_out0;
assign v_G1_1957_out0 = v_CARRY_2391_out0 || v_CARRY_2390_out0;
assign v_COUT_341_out0 = v_G1_1957_out0;
assign v_CIN_4847_out0 = v_COUT_341_out0;
assign v_RD_2902_out0 = v_CIN_4847_out0;
assign v_G1_3821_out0 = ((v_RD_2902_out0 && !v_RM_5593_out0) || (!v_RD_2902_out0) && v_RM_5593_out0);
assign v_G2_6066_out0 = v_RD_2902_out0 && v_RM_5593_out0;
assign v_CARRY_2403_out0 = v_G2_6066_out0;
assign v_S_4390_out0 = v_G1_3821_out0;
assign v_S_611_out0 = v_S_4390_out0;
assign v_G1_1963_out0 = v_CARRY_2403_out0 || v_CARRY_2402_out0;
assign v_COUT_347_out0 = v_G1_1963_out0;
assign v__2335_out0 = { v_S_605_out0,v_S_611_out0 };
assign v_CIN_4842_out0 = v_COUT_347_out0;
assign v_RD_2892_out0 = v_CIN_4842_out0;
assign v_G1_3811_out0 = ((v_RD_2892_out0 && !v_RM_5583_out0) || (!v_RD_2892_out0) && v_RM_5583_out0);
assign v_G2_6056_out0 = v_RD_2892_out0 && v_RM_5583_out0;
assign v_CARRY_2393_out0 = v_G2_6056_out0;
assign v_S_4380_out0 = v_G1_3811_out0;
assign v_S_606_out0 = v_S_4380_out0;
assign v_G1_1958_out0 = v_CARRY_2393_out0 || v_CARRY_2392_out0;
assign v_COUT_342_out0 = v_G1_1958_out0;
assign v__1244_out0 = { v__2335_out0,v_S_606_out0 };
assign v_CIN_4837_out0 = v_COUT_342_out0;
assign v_RD_2881_out0 = v_CIN_4837_out0;
assign v_G1_3800_out0 = ((v_RD_2881_out0 && !v_RM_5572_out0) || (!v_RD_2881_out0) && v_RM_5572_out0);
assign v_G2_6045_out0 = v_RD_2881_out0 && v_RM_5572_out0;
assign v_CARRY_2382_out0 = v_G2_6045_out0;
assign v_S_4369_out0 = v_G1_3800_out0;
assign v_S_601_out0 = v_S_4369_out0;
assign v_G1_1953_out0 = v_CARRY_2382_out0 || v_CARRY_2381_out0;
assign v_COUT_337_out0 = v_G1_1953_out0;
assign v__3452_out0 = { v__1244_out0,v_S_601_out0 };
assign v_CIN_4836_out0 = v_COUT_337_out0;
assign v_RD_2879_out0 = v_CIN_4836_out0;
assign v_G1_3798_out0 = ((v_RD_2879_out0 && !v_RM_5570_out0) || (!v_RD_2879_out0) && v_RM_5570_out0);
assign v_G2_6043_out0 = v_RD_2879_out0 && v_RM_5570_out0;
assign v_CARRY_2380_out0 = v_G2_6043_out0;
assign v_S_4367_out0 = v_G1_3798_out0;
assign v_S_600_out0 = v_S_4367_out0;
assign v_G1_1952_out0 = v_CARRY_2380_out0 || v_CARRY_2379_out0;
assign v_COUT_336_out0 = v_G1_1952_out0;
assign v__6662_out0 = { v__3452_out0,v_S_600_out0 };
assign v_CIN_4843_out0 = v_COUT_336_out0;
assign v_RD_2894_out0 = v_CIN_4843_out0;
assign v_G1_3813_out0 = ((v_RD_2894_out0 && !v_RM_5585_out0) || (!v_RD_2894_out0) && v_RM_5585_out0);
assign v_G2_6058_out0 = v_RD_2894_out0 && v_RM_5585_out0;
assign v_CARRY_2395_out0 = v_G2_6058_out0;
assign v_S_4382_out0 = v_G1_3813_out0;
assign v_S_607_out0 = v_S_4382_out0;
assign v_G1_1959_out0 = v_CARRY_2395_out0 || v_CARRY_2394_out0;
assign v_COUT_343_out0 = v_G1_1959_out0;
assign v__1610_out0 = { v__6662_out0,v_S_607_out0 };
assign v_CIN_4844_out0 = v_COUT_343_out0;
assign v_RD_2896_out0 = v_CIN_4844_out0;
assign v_G1_3815_out0 = ((v_RD_2896_out0 && !v_RM_5587_out0) || (!v_RD_2896_out0) && v_RM_5587_out0);
assign v_G2_6060_out0 = v_RD_2896_out0 && v_RM_5587_out0;
assign v_CARRY_2397_out0 = v_G2_6060_out0;
assign v_S_4384_out0 = v_G1_3815_out0;
assign v_S_608_out0 = v_S_4384_out0;
assign v_G1_1960_out0 = v_CARRY_2397_out0 || v_CARRY_2396_out0;
assign v_COUT_344_out0 = v_G1_1960_out0;
assign v__3507_out0 = { v__1610_out0,v_S_608_out0 };
assign v_CIN_4846_out0 = v_COUT_344_out0;
assign v_RD_2900_out0 = v_CIN_4846_out0;
assign v_G1_3819_out0 = ((v_RD_2900_out0 && !v_RM_5591_out0) || (!v_RD_2900_out0) && v_RM_5591_out0);
assign v_G2_6064_out0 = v_RD_2900_out0 && v_RM_5591_out0;
assign v_CARRY_2401_out0 = v_G2_6064_out0;
assign v_S_4388_out0 = v_G1_3819_out0;
assign v_S_610_out0 = v_S_4388_out0;
assign v_G1_1962_out0 = v_CARRY_2401_out0 || v_CARRY_2400_out0;
assign v_COUT_346_out0 = v_G1_1962_out0;
assign v__2318_out0 = { v__3507_out0,v_S_610_out0 };
assign v_CIN_4839_out0 = v_COUT_346_out0;
assign v_RD_2886_out0 = v_CIN_4839_out0;
assign v_G1_3805_out0 = ((v_RD_2886_out0 && !v_RM_5577_out0) || (!v_RD_2886_out0) && v_RM_5577_out0);
assign v_G2_6050_out0 = v_RD_2886_out0 && v_RM_5577_out0;
assign v_CARRY_2387_out0 = v_G2_6050_out0;
assign v_S_4374_out0 = v_G1_3805_out0;
assign v_S_603_out0 = v_S_4374_out0;
assign v_G1_1955_out0 = v_CARRY_2387_out0 || v_CARRY_2386_out0;
assign v_COUT_339_out0 = v_G1_1955_out0;
assign v__3400_out0 = { v__2318_out0,v_S_603_out0 };
assign v_CIN_4840_out0 = v_COUT_339_out0;
assign v_RD_2888_out0 = v_CIN_4840_out0;
assign v_G1_3807_out0 = ((v_RD_2888_out0 && !v_RM_5579_out0) || (!v_RD_2888_out0) && v_RM_5579_out0);
assign v_G2_6052_out0 = v_RD_2888_out0 && v_RM_5579_out0;
assign v_CARRY_2389_out0 = v_G2_6052_out0;
assign v_S_4376_out0 = v_G1_3807_out0;
assign v_S_604_out0 = v_S_4376_out0;
assign v_G1_1956_out0 = v_CARRY_2389_out0 || v_CARRY_2388_out0;
assign v_COUT_340_out0 = v_G1_1956_out0;
assign v__2844_out0 = { v__3400_out0,v_S_604_out0 };
assign v_CIN_4845_out0 = v_COUT_340_out0;
assign v_RD_2898_out0 = v_CIN_4845_out0;
assign v_G1_3817_out0 = ((v_RD_2898_out0 && !v_RM_5589_out0) || (!v_RD_2898_out0) && v_RM_5589_out0);
assign v_G2_6062_out0 = v_RD_2898_out0 && v_RM_5589_out0;
assign v_CARRY_2399_out0 = v_G2_6062_out0;
assign v_S_4386_out0 = v_G1_3817_out0;
assign v_S_609_out0 = v_S_4386_out0;
assign v_G1_1961_out0 = v_CARRY_2399_out0 || v_CARRY_2398_out0;
assign v_COUT_345_out0 = v_G1_1961_out0;
assign v__988_out0 = { v__2844_out0,v_S_609_out0 };
assign v_CIN_4833_out0 = v_COUT_345_out0;
assign v_RD_2873_out0 = v_CIN_4833_out0;
assign v_G1_3792_out0 = ((v_RD_2873_out0 && !v_RM_5564_out0) || (!v_RD_2873_out0) && v_RM_5564_out0);
assign v_G2_6037_out0 = v_RD_2873_out0 && v_RM_5564_out0;
assign v_CARRY_2374_out0 = v_G2_6037_out0;
assign v_S_4361_out0 = v_G1_3792_out0;
assign v_S_597_out0 = v_S_4361_out0;
assign v_G1_1949_out0 = v_CARRY_2374_out0 || v_CARRY_2373_out0;
assign v_COUT_333_out0 = v_G1_1949_out0;
assign v__1364_out0 = { v__988_out0,v_S_597_out0 };
assign v_CIN_4838_out0 = v_COUT_333_out0;
assign v_RD_2883_out0 = v_CIN_4838_out0;
assign v_G1_3802_out0 = ((v_RD_2883_out0 && !v_RM_5574_out0) || (!v_RD_2883_out0) && v_RM_5574_out0);
assign v_G2_6047_out0 = v_RD_2883_out0 && v_RM_5574_out0;
assign v_CARRY_2384_out0 = v_G2_6047_out0;
assign v_S_4371_out0 = v_G1_3802_out0;
assign v_S_602_out0 = v_S_4371_out0;
assign v_G1_1954_out0 = v_CARRY_2384_out0 || v_CARRY_2383_out0;
assign v_COUT_338_out0 = v_G1_1954_out0;
assign v__891_out0 = { v__1364_out0,v_S_602_out0 };
assign v_CIN_4834_out0 = v_COUT_338_out0;
assign v_RD_2875_out0 = v_CIN_4834_out0;
assign v_G1_3794_out0 = ((v_RD_2875_out0 && !v_RM_5566_out0) || (!v_RD_2875_out0) && v_RM_5566_out0);
assign v_G2_6039_out0 = v_RD_2875_out0 && v_RM_5566_out0;
assign v_CARRY_2376_out0 = v_G2_6039_out0;
assign v_S_4363_out0 = v_G1_3794_out0;
assign v_S_598_out0 = v_S_4363_out0;
assign v_G1_1950_out0 = v_CARRY_2376_out0 || v_CARRY_2375_out0;
assign v_COUT_334_out0 = v_G1_1950_out0;
assign v__2220_out0 = { v__891_out0,v_S_598_out0 };
assign v_RM_1632_out0 = v_COUT_334_out0;
assign v_RM_5567_out0 = v_RM_1632_out0;
assign v_G1_3795_out0 = ((v_RD_2876_out0 && !v_RM_5567_out0) || (!v_RD_2876_out0) && v_RM_5567_out0);
assign v_G2_6040_out0 = v_RD_2876_out0 && v_RM_5567_out0;
assign v_CARRY_2377_out0 = v_G2_6040_out0;
assign v_S_4364_out0 = v_G1_3795_out0;
assign v_RM_5568_out0 = v_S_4364_out0;
assign v_G1_3796_out0 = ((v_RD_2877_out0 && !v_RM_5568_out0) || (!v_RD_2877_out0) && v_RM_5568_out0);
assign v_G2_6041_out0 = v_RD_2877_out0 && v_RM_5568_out0;
assign v_CARRY_2378_out0 = v_G2_6041_out0;
assign v_S_4365_out0 = v_G1_3796_out0;
assign v_S_599_out0 = v_S_4365_out0;
assign v_G1_1951_out0 = v_CARRY_2378_out0 || v_CARRY_2377_out0;
assign v_COUT_335_out0 = v_G1_1951_out0;
assign v__5243_out0 = { v__2220_out0,v_S_599_out0 };
assign v__5386_out0 = { v__5243_out0,v_COUT_335_out0 };
assign v_COUT_5371_out0 = v__5386_out0;
assign v_CIN_1157_out0 = v_COUT_5371_out0;
assign v__239_out0 = v_CIN_1157_out0[8:8];
assign v__877_out0 = v_CIN_1157_out0[6:6];
assign v__1060_out0 = v_CIN_1157_out0[3:3];
assign v__1079_out0 = v_CIN_1157_out0[15:15];
assign v__1230_out0 = v_CIN_1157_out0[0:0];
assign v__1498_out0 = v_CIN_1157_out0[9:9];
assign v__1514_out0 = v_CIN_1157_out0[2:2];
assign v__1540_out0 = v_CIN_1157_out0[7:7];
assign v__1873_out0 = v_CIN_1157_out0[1:1];
assign v__1891_out0 = v_CIN_1157_out0[10:10];
assign v__3350_out0 = v_CIN_1157_out0[11:11];
assign v__3766_out0 = v_CIN_1157_out0[12:12];
assign v__4292_out0 = v_CIN_1157_out0[13:13];
assign v__4325_out0 = v_CIN_1157_out0[14:14];
assign v__5286_out0 = v_CIN_1157_out0[5:5];
assign v__6634_out0 = v_CIN_1157_out0[4:4];
assign v_RM_1779_out0 = v__3766_out0;
assign v_RM_1780_out0 = v__4325_out0;
assign v_RM_1782_out0 = v__5286_out0;
assign v_RM_1783_out0 = v__6634_out0;
assign v_RM_1784_out0 = v__4292_out0;
assign v_RM_1785_out0 = v__1498_out0;
assign v_RM_1786_out0 = v__1891_out0;
assign v_RM_1787_out0 = v__1873_out0;
assign v_RM_1788_out0 = v__1060_out0;
assign v_RM_1789_out0 = v__877_out0;
assign v_RM_1790_out0 = v__1540_out0;
assign v_RM_1791_out0 = v__3350_out0;
assign v_RM_1792_out0 = v__239_out0;
assign v_RM_1793_out0 = v__1514_out0;
assign v_CIN_4984_out0 = v__1079_out0;
assign v_RM_5884_out0 = v__1230_out0;
assign v_RD_3186_out0 = v_CIN_4984_out0;
assign v_G1_4112_out0 = ((v_RD_3193_out0 && !v_RM_5884_out0) || (!v_RD_3193_out0) && v_RM_5884_out0);
assign v_RM_5872_out0 = v_RM_1779_out0;
assign v_RM_5874_out0 = v_RM_1780_out0;
assign v_RM_5878_out0 = v_RM_1782_out0;
assign v_RM_5880_out0 = v_RM_1783_out0;
assign v_RM_5882_out0 = v_RM_1784_out0;
assign v_RM_5885_out0 = v_RM_1785_out0;
assign v_RM_5887_out0 = v_RM_1786_out0;
assign v_RM_5889_out0 = v_RM_1787_out0;
assign v_RM_5891_out0 = v_RM_1788_out0;
assign v_RM_5893_out0 = v_RM_1789_out0;
assign v_RM_5895_out0 = v_RM_1790_out0;
assign v_RM_5897_out0 = v_RM_1791_out0;
assign v_RM_5899_out0 = v_RM_1792_out0;
assign v_RM_5901_out0 = v_RM_1793_out0;
assign v_G2_6357_out0 = v_RD_3193_out0 && v_RM_5884_out0;
assign v_CARRY_2694_out0 = v_G2_6357_out0;
assign v_G1_4100_out0 = ((v_RD_3181_out0 && !v_RM_5872_out0) || (!v_RD_3181_out0) && v_RM_5872_out0);
assign v_G1_4102_out0 = ((v_RD_3183_out0 && !v_RM_5874_out0) || (!v_RD_3183_out0) && v_RM_5874_out0);
assign v_G1_4106_out0 = ((v_RD_3187_out0 && !v_RM_5878_out0) || (!v_RD_3187_out0) && v_RM_5878_out0);
assign v_G1_4108_out0 = ((v_RD_3189_out0 && !v_RM_5880_out0) || (!v_RD_3189_out0) && v_RM_5880_out0);
assign v_G1_4110_out0 = ((v_RD_3191_out0 && !v_RM_5882_out0) || (!v_RD_3191_out0) && v_RM_5882_out0);
assign v_G1_4113_out0 = ((v_RD_3194_out0 && !v_RM_5885_out0) || (!v_RD_3194_out0) && v_RM_5885_out0);
assign v_G1_4115_out0 = ((v_RD_3196_out0 && !v_RM_5887_out0) || (!v_RD_3196_out0) && v_RM_5887_out0);
assign v_G1_4117_out0 = ((v_RD_3198_out0 && !v_RM_5889_out0) || (!v_RD_3198_out0) && v_RM_5889_out0);
assign v_G1_4119_out0 = ((v_RD_3200_out0 && !v_RM_5891_out0) || (!v_RD_3200_out0) && v_RM_5891_out0);
assign v_G1_4121_out0 = ((v_RD_3202_out0 && !v_RM_5893_out0) || (!v_RD_3202_out0) && v_RM_5893_out0);
assign v_G1_4123_out0 = ((v_RD_3204_out0 && !v_RM_5895_out0) || (!v_RD_3204_out0) && v_RM_5895_out0);
assign v_G1_4125_out0 = ((v_RD_3206_out0 && !v_RM_5897_out0) || (!v_RD_3206_out0) && v_RM_5897_out0);
assign v_G1_4127_out0 = ((v_RD_3208_out0 && !v_RM_5899_out0) || (!v_RD_3208_out0) && v_RM_5899_out0);
assign v_G1_4129_out0 = ((v_RD_3210_out0 && !v_RM_5901_out0) || (!v_RD_3210_out0) && v_RM_5901_out0);
assign v_S_4681_out0 = v_G1_4112_out0;
assign v_G2_6345_out0 = v_RD_3181_out0 && v_RM_5872_out0;
assign v_G2_6347_out0 = v_RD_3183_out0 && v_RM_5874_out0;
assign v_G2_6351_out0 = v_RD_3187_out0 && v_RM_5878_out0;
assign v_G2_6353_out0 = v_RD_3189_out0 && v_RM_5880_out0;
assign v_G2_6355_out0 = v_RD_3191_out0 && v_RM_5882_out0;
assign v_G2_6358_out0 = v_RD_3194_out0 && v_RM_5885_out0;
assign v_G2_6360_out0 = v_RD_3196_out0 && v_RM_5887_out0;
assign v_G2_6362_out0 = v_RD_3198_out0 && v_RM_5889_out0;
assign v_G2_6364_out0 = v_RD_3200_out0 && v_RM_5891_out0;
assign v_G2_6366_out0 = v_RD_3202_out0 && v_RM_5893_out0;
assign v_G2_6368_out0 = v_RD_3204_out0 && v_RM_5895_out0;
assign v_G2_6370_out0 = v_RD_3206_out0 && v_RM_5897_out0;
assign v_G2_6372_out0 = v_RD_3208_out0 && v_RM_5899_out0;
assign v_G2_6374_out0 = v_RD_3210_out0 && v_RM_5901_out0;
assign v_S_2288_out0 = v_S_4681_out0;
assign v_CARRY_2682_out0 = v_G2_6345_out0;
assign v_CARRY_2684_out0 = v_G2_6347_out0;
assign v_CARRY_2688_out0 = v_G2_6351_out0;
assign v_CARRY_2690_out0 = v_G2_6353_out0;
assign v_CARRY_2692_out0 = v_G2_6355_out0;
assign v_CARRY_2695_out0 = v_G2_6358_out0;
assign v_CARRY_2697_out0 = v_G2_6360_out0;
assign v_CARRY_2699_out0 = v_G2_6362_out0;
assign v_CARRY_2701_out0 = v_G2_6364_out0;
assign v_CARRY_2703_out0 = v_G2_6366_out0;
assign v_CARRY_2705_out0 = v_G2_6368_out0;
assign v_CARRY_2707_out0 = v_G2_6370_out0;
assign v_CARRY_2709_out0 = v_G2_6372_out0;
assign v_CARRY_2711_out0 = v_G2_6374_out0;
assign v_S_4669_out0 = v_G1_4100_out0;
assign v_S_4671_out0 = v_G1_4102_out0;
assign v_S_4675_out0 = v_G1_4106_out0;
assign v_S_4677_out0 = v_G1_4108_out0;
assign v_S_4679_out0 = v_G1_4110_out0;
assign v_S_4682_out0 = v_G1_4113_out0;
assign v_S_4684_out0 = v_G1_4115_out0;
assign v_S_4686_out0 = v_G1_4117_out0;
assign v_S_4688_out0 = v_G1_4119_out0;
assign v_S_4690_out0 = v_G1_4121_out0;
assign v_S_4692_out0 = v_G1_4123_out0;
assign v_S_4694_out0 = v_G1_4125_out0;
assign v_S_4696_out0 = v_G1_4127_out0;
assign v_S_4698_out0 = v_G1_4129_out0;
assign v_CIN_4990_out0 = v_CARRY_2694_out0;
assign v__30_out0 = { v__1166_out0,v_S_2288_out0 };
assign v_RD_3199_out0 = v_CIN_4990_out0;
assign v_RM_5873_out0 = v_S_4669_out0;
assign v_RM_5875_out0 = v_S_4671_out0;
assign v_RM_5879_out0 = v_S_4675_out0;
assign v_RM_5881_out0 = v_S_4677_out0;
assign v_RM_5883_out0 = v_S_4679_out0;
assign v_RM_5886_out0 = v_S_4682_out0;
assign v_RM_5888_out0 = v_S_4684_out0;
assign v_RM_5890_out0 = v_S_4686_out0;
assign v_RM_5892_out0 = v_S_4688_out0;
assign v_RM_5894_out0 = v_S_4690_out0;
assign v_RM_5896_out0 = v_S_4692_out0;
assign v_RM_5898_out0 = v_S_4694_out0;
assign v_RM_5900_out0 = v_S_4696_out0;
assign v_RM_5902_out0 = v_S_4698_out0;
assign v_G1_4118_out0 = ((v_RD_3199_out0 && !v_RM_5890_out0) || (!v_RD_3199_out0) && v_RM_5890_out0);
assign v_G2_6363_out0 = v_RD_3199_out0 && v_RM_5890_out0;
assign v_CARRY_2700_out0 = v_G2_6363_out0;
assign v_S_4687_out0 = v_G1_4118_out0;
assign v_S_754_out0 = v_S_4687_out0;
assign v_G1_2106_out0 = v_CARRY_2700_out0 || v_CARRY_2699_out0;
assign v_COUT_490_out0 = v_G1_2106_out0;
assign v_CIN_4996_out0 = v_COUT_490_out0;
assign v_RD_3211_out0 = v_CIN_4996_out0;
assign v_G1_4130_out0 = ((v_RD_3211_out0 && !v_RM_5902_out0) || (!v_RD_3211_out0) && v_RM_5902_out0);
assign v_G2_6375_out0 = v_RD_3211_out0 && v_RM_5902_out0;
assign v_CARRY_2712_out0 = v_G2_6375_out0;
assign v_S_4699_out0 = v_G1_4130_out0;
assign v_S_760_out0 = v_S_4699_out0;
assign v_G1_2112_out0 = v_CARRY_2712_out0 || v_CARRY_2711_out0;
assign v_COUT_496_out0 = v_G1_2112_out0;
assign v__2345_out0 = { v_S_754_out0,v_S_760_out0 };
assign v_CIN_4991_out0 = v_COUT_496_out0;
assign v_RD_3201_out0 = v_CIN_4991_out0;
assign v_G1_4120_out0 = ((v_RD_3201_out0 && !v_RM_5892_out0) || (!v_RD_3201_out0) && v_RM_5892_out0);
assign v_G2_6365_out0 = v_RD_3201_out0 && v_RM_5892_out0;
assign v_CARRY_2702_out0 = v_G2_6365_out0;
assign v_S_4689_out0 = v_G1_4120_out0;
assign v_S_755_out0 = v_S_4689_out0;
assign v_G1_2107_out0 = v_CARRY_2702_out0 || v_CARRY_2701_out0;
assign v_COUT_491_out0 = v_G1_2107_out0;
assign v__1254_out0 = { v__2345_out0,v_S_755_out0 };
assign v_CIN_4986_out0 = v_COUT_491_out0;
assign v_RD_3190_out0 = v_CIN_4986_out0;
assign v_G1_4109_out0 = ((v_RD_3190_out0 && !v_RM_5881_out0) || (!v_RD_3190_out0) && v_RM_5881_out0);
assign v_G2_6354_out0 = v_RD_3190_out0 && v_RM_5881_out0;
assign v_CARRY_2691_out0 = v_G2_6354_out0;
assign v_S_4678_out0 = v_G1_4109_out0;
assign v_S_750_out0 = v_S_4678_out0;
assign v_G1_2102_out0 = v_CARRY_2691_out0 || v_CARRY_2690_out0;
assign v_COUT_486_out0 = v_G1_2102_out0;
assign v__3462_out0 = { v__1254_out0,v_S_750_out0 };
assign v_CIN_4985_out0 = v_COUT_486_out0;
assign v_RD_3188_out0 = v_CIN_4985_out0;
assign v_G1_4107_out0 = ((v_RD_3188_out0 && !v_RM_5879_out0) || (!v_RD_3188_out0) && v_RM_5879_out0);
assign v_G2_6352_out0 = v_RD_3188_out0 && v_RM_5879_out0;
assign v_CARRY_2689_out0 = v_G2_6352_out0;
assign v_S_4676_out0 = v_G1_4107_out0;
assign v_S_749_out0 = v_S_4676_out0;
assign v_G1_2101_out0 = v_CARRY_2689_out0 || v_CARRY_2688_out0;
assign v_COUT_485_out0 = v_G1_2101_out0;
assign v__6672_out0 = { v__3462_out0,v_S_749_out0 };
assign v_CIN_4992_out0 = v_COUT_485_out0;
assign v_RD_3203_out0 = v_CIN_4992_out0;
assign v_G1_4122_out0 = ((v_RD_3203_out0 && !v_RM_5894_out0) || (!v_RD_3203_out0) && v_RM_5894_out0);
assign v_G2_6367_out0 = v_RD_3203_out0 && v_RM_5894_out0;
assign v_CARRY_2704_out0 = v_G2_6367_out0;
assign v_S_4691_out0 = v_G1_4122_out0;
assign v_S_756_out0 = v_S_4691_out0;
assign v_G1_2108_out0 = v_CARRY_2704_out0 || v_CARRY_2703_out0;
assign v_COUT_492_out0 = v_G1_2108_out0;
assign v__1620_out0 = { v__6672_out0,v_S_756_out0 };
assign v_CIN_4993_out0 = v_COUT_492_out0;
assign v_RD_3205_out0 = v_CIN_4993_out0;
assign v_G1_4124_out0 = ((v_RD_3205_out0 && !v_RM_5896_out0) || (!v_RD_3205_out0) && v_RM_5896_out0);
assign v_G2_6369_out0 = v_RD_3205_out0 && v_RM_5896_out0;
assign v_CARRY_2706_out0 = v_G2_6369_out0;
assign v_S_4693_out0 = v_G1_4124_out0;
assign v_S_757_out0 = v_S_4693_out0;
assign v_G1_2109_out0 = v_CARRY_2706_out0 || v_CARRY_2705_out0;
assign v_COUT_493_out0 = v_G1_2109_out0;
assign v__3517_out0 = { v__1620_out0,v_S_757_out0 };
assign v_CIN_4995_out0 = v_COUT_493_out0;
assign v_RD_3209_out0 = v_CIN_4995_out0;
assign v_G1_4128_out0 = ((v_RD_3209_out0 && !v_RM_5900_out0) || (!v_RD_3209_out0) && v_RM_5900_out0);
assign v_G2_6373_out0 = v_RD_3209_out0 && v_RM_5900_out0;
assign v_CARRY_2710_out0 = v_G2_6373_out0;
assign v_S_4697_out0 = v_G1_4128_out0;
assign v_S_759_out0 = v_S_4697_out0;
assign v_G1_2111_out0 = v_CARRY_2710_out0 || v_CARRY_2709_out0;
assign v_COUT_495_out0 = v_G1_2111_out0;
assign v__2328_out0 = { v__3517_out0,v_S_759_out0 };
assign v_CIN_4988_out0 = v_COUT_495_out0;
assign v_RD_3195_out0 = v_CIN_4988_out0;
assign v_G1_4114_out0 = ((v_RD_3195_out0 && !v_RM_5886_out0) || (!v_RD_3195_out0) && v_RM_5886_out0);
assign v_G2_6359_out0 = v_RD_3195_out0 && v_RM_5886_out0;
assign v_CARRY_2696_out0 = v_G2_6359_out0;
assign v_S_4683_out0 = v_G1_4114_out0;
assign v_S_752_out0 = v_S_4683_out0;
assign v_G1_2104_out0 = v_CARRY_2696_out0 || v_CARRY_2695_out0;
assign v_COUT_488_out0 = v_G1_2104_out0;
assign v__3410_out0 = { v__2328_out0,v_S_752_out0 };
assign v_CIN_4989_out0 = v_COUT_488_out0;
assign v_RD_3197_out0 = v_CIN_4989_out0;
assign v_G1_4116_out0 = ((v_RD_3197_out0 && !v_RM_5888_out0) || (!v_RD_3197_out0) && v_RM_5888_out0);
assign v_G2_6361_out0 = v_RD_3197_out0 && v_RM_5888_out0;
assign v_CARRY_2698_out0 = v_G2_6361_out0;
assign v_S_4685_out0 = v_G1_4116_out0;
assign v_S_753_out0 = v_S_4685_out0;
assign v_G1_2105_out0 = v_CARRY_2698_out0 || v_CARRY_2697_out0;
assign v_COUT_489_out0 = v_G1_2105_out0;
assign v__2854_out0 = { v__3410_out0,v_S_753_out0 };
assign v_CIN_4994_out0 = v_COUT_489_out0;
assign v_RD_3207_out0 = v_CIN_4994_out0;
assign v_G1_4126_out0 = ((v_RD_3207_out0 && !v_RM_5898_out0) || (!v_RD_3207_out0) && v_RM_5898_out0);
assign v_G2_6371_out0 = v_RD_3207_out0 && v_RM_5898_out0;
assign v_CARRY_2708_out0 = v_G2_6371_out0;
assign v_S_4695_out0 = v_G1_4126_out0;
assign v_S_758_out0 = v_S_4695_out0;
assign v_G1_2110_out0 = v_CARRY_2708_out0 || v_CARRY_2707_out0;
assign v_COUT_494_out0 = v_G1_2110_out0;
assign v__998_out0 = { v__2854_out0,v_S_758_out0 };
assign v_CIN_4982_out0 = v_COUT_494_out0;
assign v_RD_3182_out0 = v_CIN_4982_out0;
assign v_G1_4101_out0 = ((v_RD_3182_out0 && !v_RM_5873_out0) || (!v_RD_3182_out0) && v_RM_5873_out0);
assign v_G2_6346_out0 = v_RD_3182_out0 && v_RM_5873_out0;
assign v_CARRY_2683_out0 = v_G2_6346_out0;
assign v_S_4670_out0 = v_G1_4101_out0;
assign v_S_746_out0 = v_S_4670_out0;
assign v_G1_2098_out0 = v_CARRY_2683_out0 || v_CARRY_2682_out0;
assign v_COUT_482_out0 = v_G1_2098_out0;
assign v__1374_out0 = { v__998_out0,v_S_746_out0 };
assign v_CIN_4987_out0 = v_COUT_482_out0;
assign v_RD_3192_out0 = v_CIN_4987_out0;
assign v_G1_4111_out0 = ((v_RD_3192_out0 && !v_RM_5883_out0) || (!v_RD_3192_out0) && v_RM_5883_out0);
assign v_G2_6356_out0 = v_RD_3192_out0 && v_RM_5883_out0;
assign v_CARRY_2693_out0 = v_G2_6356_out0;
assign v_S_4680_out0 = v_G1_4111_out0;
assign v_S_751_out0 = v_S_4680_out0;
assign v_G1_2103_out0 = v_CARRY_2693_out0 || v_CARRY_2692_out0;
assign v_COUT_487_out0 = v_G1_2103_out0;
assign v__901_out0 = { v__1374_out0,v_S_751_out0 };
assign v_CIN_4983_out0 = v_COUT_487_out0;
assign v_RD_3184_out0 = v_CIN_4983_out0;
assign v_G1_4103_out0 = ((v_RD_3184_out0 && !v_RM_5875_out0) || (!v_RD_3184_out0) && v_RM_5875_out0);
assign v_G2_6348_out0 = v_RD_3184_out0 && v_RM_5875_out0;
assign v_CARRY_2685_out0 = v_G2_6348_out0;
assign v_S_4672_out0 = v_G1_4103_out0;
assign v_S_747_out0 = v_S_4672_out0;
assign v_G1_2099_out0 = v_CARRY_2685_out0 || v_CARRY_2684_out0;
assign v_COUT_483_out0 = v_G1_2099_out0;
assign v__2230_out0 = { v__901_out0,v_S_747_out0 };
assign v_RM_1781_out0 = v_COUT_483_out0;
assign v_RM_5876_out0 = v_RM_1781_out0;
assign v_G1_4104_out0 = ((v_RD_3185_out0 && !v_RM_5876_out0) || (!v_RD_3185_out0) && v_RM_5876_out0);
assign v_G2_6349_out0 = v_RD_3185_out0 && v_RM_5876_out0;
assign v_CARRY_2686_out0 = v_G2_6349_out0;
assign v_S_4673_out0 = v_G1_4104_out0;
assign v_RM_5877_out0 = v_S_4673_out0;
assign v_G1_4105_out0 = ((v_RD_3186_out0 && !v_RM_5877_out0) || (!v_RD_3186_out0) && v_RM_5877_out0);
assign v_G2_6350_out0 = v_RD_3186_out0 && v_RM_5877_out0;
assign v_CARRY_2687_out0 = v_G2_6350_out0;
assign v_S_4674_out0 = v_G1_4105_out0;
assign v_S_748_out0 = v_S_4674_out0;
assign v_G1_2100_out0 = v_CARRY_2687_out0 || v_CARRY_2686_out0;
assign v_COUT_484_out0 = v_G1_2100_out0;
assign v__5253_out0 = { v__2230_out0,v_S_748_out0 };
assign v__5396_out0 = { v__5253_out0,v_COUT_484_out0 };
assign v_COUT_5381_out0 = v__5396_out0;
assign v_CIN_1160_out0 = v_COUT_5381_out0;
assign v__242_out0 = v_CIN_1160_out0[8:8];
assign v__880_out0 = v_CIN_1160_out0[6:6];
assign v__1063_out0 = v_CIN_1160_out0[3:3];
assign v__1082_out0 = v_CIN_1160_out0[15:15];
assign v__1233_out0 = v_CIN_1160_out0[0:0];
assign v__1501_out0 = v_CIN_1160_out0[9:9];
assign v__1517_out0 = v_CIN_1160_out0[2:2];
assign v__1543_out0 = v_CIN_1160_out0[7:7];
assign v__1876_out0 = v_CIN_1160_out0[1:1];
assign v__1894_out0 = v_CIN_1160_out0[10:10];
assign v__3353_out0 = v_CIN_1160_out0[11:11];
assign v__3769_out0 = v_CIN_1160_out0[12:12];
assign v__4295_out0 = v_CIN_1160_out0[13:13];
assign v__4328_out0 = v_CIN_1160_out0[14:14];
assign v__5289_out0 = v_CIN_1160_out0[5:5];
assign v__6637_out0 = v_CIN_1160_out0[4:4];
assign v_RM_1824_out0 = v__3769_out0;
assign v_RM_1825_out0 = v__4328_out0;
assign v_RM_1827_out0 = v__5289_out0;
assign v_RM_1828_out0 = v__6637_out0;
assign v_RM_1829_out0 = v__4295_out0;
assign v_RM_1830_out0 = v__1501_out0;
assign v_RM_1831_out0 = v__1894_out0;
assign v_RM_1832_out0 = v__1876_out0;
assign v_RM_1833_out0 = v__1063_out0;
assign v_RM_1834_out0 = v__880_out0;
assign v_RM_1835_out0 = v__1543_out0;
assign v_RM_1836_out0 = v__3353_out0;
assign v_RM_1837_out0 = v__242_out0;
assign v_RM_1838_out0 = v__1517_out0;
assign v_CIN_5029_out0 = v__1082_out0;
assign v_RM_5977_out0 = v__1233_out0;
assign v_RD_3279_out0 = v_CIN_5029_out0;
assign v_G1_4205_out0 = ((v_RD_3286_out0 && !v_RM_5977_out0) || (!v_RD_3286_out0) && v_RM_5977_out0);
assign v_RM_5965_out0 = v_RM_1824_out0;
assign v_RM_5967_out0 = v_RM_1825_out0;
assign v_RM_5971_out0 = v_RM_1827_out0;
assign v_RM_5973_out0 = v_RM_1828_out0;
assign v_RM_5975_out0 = v_RM_1829_out0;
assign v_RM_5978_out0 = v_RM_1830_out0;
assign v_RM_5980_out0 = v_RM_1831_out0;
assign v_RM_5982_out0 = v_RM_1832_out0;
assign v_RM_5984_out0 = v_RM_1833_out0;
assign v_RM_5986_out0 = v_RM_1834_out0;
assign v_RM_5988_out0 = v_RM_1835_out0;
assign v_RM_5990_out0 = v_RM_1836_out0;
assign v_RM_5992_out0 = v_RM_1837_out0;
assign v_RM_5994_out0 = v_RM_1838_out0;
assign v_G2_6450_out0 = v_RD_3286_out0 && v_RM_5977_out0;
assign v_CARRY_2787_out0 = v_G2_6450_out0;
assign v_G1_4193_out0 = ((v_RD_3274_out0 && !v_RM_5965_out0) || (!v_RD_3274_out0) && v_RM_5965_out0);
assign v_G1_4195_out0 = ((v_RD_3276_out0 && !v_RM_5967_out0) || (!v_RD_3276_out0) && v_RM_5967_out0);
assign v_G1_4199_out0 = ((v_RD_3280_out0 && !v_RM_5971_out0) || (!v_RD_3280_out0) && v_RM_5971_out0);
assign v_G1_4201_out0 = ((v_RD_3282_out0 && !v_RM_5973_out0) || (!v_RD_3282_out0) && v_RM_5973_out0);
assign v_G1_4203_out0 = ((v_RD_3284_out0 && !v_RM_5975_out0) || (!v_RD_3284_out0) && v_RM_5975_out0);
assign v_G1_4206_out0 = ((v_RD_3287_out0 && !v_RM_5978_out0) || (!v_RD_3287_out0) && v_RM_5978_out0);
assign v_G1_4208_out0 = ((v_RD_3289_out0 && !v_RM_5980_out0) || (!v_RD_3289_out0) && v_RM_5980_out0);
assign v_G1_4210_out0 = ((v_RD_3291_out0 && !v_RM_5982_out0) || (!v_RD_3291_out0) && v_RM_5982_out0);
assign v_G1_4212_out0 = ((v_RD_3293_out0 && !v_RM_5984_out0) || (!v_RD_3293_out0) && v_RM_5984_out0);
assign v_G1_4214_out0 = ((v_RD_3295_out0 && !v_RM_5986_out0) || (!v_RD_3295_out0) && v_RM_5986_out0);
assign v_G1_4216_out0 = ((v_RD_3297_out0 && !v_RM_5988_out0) || (!v_RD_3297_out0) && v_RM_5988_out0);
assign v_G1_4218_out0 = ((v_RD_3299_out0 && !v_RM_5990_out0) || (!v_RD_3299_out0) && v_RM_5990_out0);
assign v_G1_4220_out0 = ((v_RD_3301_out0 && !v_RM_5992_out0) || (!v_RD_3301_out0) && v_RM_5992_out0);
assign v_G1_4222_out0 = ((v_RD_3303_out0 && !v_RM_5994_out0) || (!v_RD_3303_out0) && v_RM_5994_out0);
assign v_S_4774_out0 = v_G1_4205_out0;
assign v_G2_6438_out0 = v_RD_3274_out0 && v_RM_5965_out0;
assign v_G2_6440_out0 = v_RD_3276_out0 && v_RM_5967_out0;
assign v_G2_6444_out0 = v_RD_3280_out0 && v_RM_5971_out0;
assign v_G2_6446_out0 = v_RD_3282_out0 && v_RM_5973_out0;
assign v_G2_6448_out0 = v_RD_3284_out0 && v_RM_5975_out0;
assign v_G2_6451_out0 = v_RD_3287_out0 && v_RM_5978_out0;
assign v_G2_6453_out0 = v_RD_3289_out0 && v_RM_5980_out0;
assign v_G2_6455_out0 = v_RD_3291_out0 && v_RM_5982_out0;
assign v_G2_6457_out0 = v_RD_3293_out0 && v_RM_5984_out0;
assign v_G2_6459_out0 = v_RD_3295_out0 && v_RM_5986_out0;
assign v_G2_6461_out0 = v_RD_3297_out0 && v_RM_5988_out0;
assign v_G2_6463_out0 = v_RD_3299_out0 && v_RM_5990_out0;
assign v_G2_6465_out0 = v_RD_3301_out0 && v_RM_5992_out0;
assign v_G2_6467_out0 = v_RD_3303_out0 && v_RM_5994_out0;
assign v_S_2291_out0 = v_S_4774_out0;
assign v_CARRY_2775_out0 = v_G2_6438_out0;
assign v_CARRY_2777_out0 = v_G2_6440_out0;
assign v_CARRY_2781_out0 = v_G2_6444_out0;
assign v_CARRY_2783_out0 = v_G2_6446_out0;
assign v_CARRY_2785_out0 = v_G2_6448_out0;
assign v_CARRY_2788_out0 = v_G2_6451_out0;
assign v_CARRY_2790_out0 = v_G2_6453_out0;
assign v_CARRY_2792_out0 = v_G2_6455_out0;
assign v_CARRY_2794_out0 = v_G2_6457_out0;
assign v_CARRY_2796_out0 = v_G2_6459_out0;
assign v_CARRY_2798_out0 = v_G2_6461_out0;
assign v_CARRY_2800_out0 = v_G2_6463_out0;
assign v_CARRY_2802_out0 = v_G2_6465_out0;
assign v_CARRY_2804_out0 = v_G2_6467_out0;
assign v_S_4762_out0 = v_G1_4193_out0;
assign v_S_4764_out0 = v_G1_4195_out0;
assign v_S_4768_out0 = v_G1_4199_out0;
assign v_S_4770_out0 = v_G1_4201_out0;
assign v_S_4772_out0 = v_G1_4203_out0;
assign v_S_4775_out0 = v_G1_4206_out0;
assign v_S_4777_out0 = v_G1_4208_out0;
assign v_S_4779_out0 = v_G1_4210_out0;
assign v_S_4781_out0 = v_G1_4212_out0;
assign v_S_4783_out0 = v_G1_4214_out0;
assign v_S_4785_out0 = v_G1_4216_out0;
assign v_S_4787_out0 = v_G1_4218_out0;
assign v_S_4789_out0 = v_G1_4220_out0;
assign v_S_4791_out0 = v_G1_4222_out0;
assign v_CIN_5035_out0 = v_CARRY_2787_out0;
assign v__330_out0 = { v__30_out0,v_S_2291_out0 };
assign v_RD_3292_out0 = v_CIN_5035_out0;
assign v_RM_5966_out0 = v_S_4762_out0;
assign v_RM_5968_out0 = v_S_4764_out0;
assign v_RM_5972_out0 = v_S_4768_out0;
assign v_RM_5974_out0 = v_S_4770_out0;
assign v_RM_5976_out0 = v_S_4772_out0;
assign v_RM_5979_out0 = v_S_4775_out0;
assign v_RM_5981_out0 = v_S_4777_out0;
assign v_RM_5983_out0 = v_S_4779_out0;
assign v_RM_5985_out0 = v_S_4781_out0;
assign v_RM_5987_out0 = v_S_4783_out0;
assign v_RM_5989_out0 = v_S_4785_out0;
assign v_RM_5991_out0 = v_S_4787_out0;
assign v_RM_5993_out0 = v_S_4789_out0;
assign v_RM_5995_out0 = v_S_4791_out0;
assign v_G1_4211_out0 = ((v_RD_3292_out0 && !v_RM_5983_out0) || (!v_RD_3292_out0) && v_RM_5983_out0);
assign v_G2_6456_out0 = v_RD_3292_out0 && v_RM_5983_out0;
assign v_CARRY_2793_out0 = v_G2_6456_out0;
assign v_S_4780_out0 = v_G1_4211_out0;
assign v_S_799_out0 = v_S_4780_out0;
assign v_G1_2151_out0 = v_CARRY_2793_out0 || v_CARRY_2792_out0;
assign v_COUT_535_out0 = v_G1_2151_out0;
assign v_CIN_5041_out0 = v_COUT_535_out0;
assign v_RD_3304_out0 = v_CIN_5041_out0;
assign v_G1_4223_out0 = ((v_RD_3304_out0 && !v_RM_5995_out0) || (!v_RD_3304_out0) && v_RM_5995_out0);
assign v_G2_6468_out0 = v_RD_3304_out0 && v_RM_5995_out0;
assign v_CARRY_2805_out0 = v_G2_6468_out0;
assign v_S_4792_out0 = v_G1_4223_out0;
assign v_S_805_out0 = v_S_4792_out0;
assign v_G1_2157_out0 = v_CARRY_2805_out0 || v_CARRY_2804_out0;
assign v_COUT_541_out0 = v_G1_2157_out0;
assign v__2348_out0 = { v_S_799_out0,v_S_805_out0 };
assign v_CIN_5036_out0 = v_COUT_541_out0;
assign v_RD_3294_out0 = v_CIN_5036_out0;
assign v_G1_4213_out0 = ((v_RD_3294_out0 && !v_RM_5985_out0) || (!v_RD_3294_out0) && v_RM_5985_out0);
assign v_G2_6458_out0 = v_RD_3294_out0 && v_RM_5985_out0;
assign v_CARRY_2795_out0 = v_G2_6458_out0;
assign v_S_4782_out0 = v_G1_4213_out0;
assign v_S_800_out0 = v_S_4782_out0;
assign v_G1_2152_out0 = v_CARRY_2795_out0 || v_CARRY_2794_out0;
assign v_COUT_536_out0 = v_G1_2152_out0;
assign v__1257_out0 = { v__2348_out0,v_S_800_out0 };
assign v_CIN_5031_out0 = v_COUT_536_out0;
assign v_RD_3283_out0 = v_CIN_5031_out0;
assign v_G1_4202_out0 = ((v_RD_3283_out0 && !v_RM_5974_out0) || (!v_RD_3283_out0) && v_RM_5974_out0);
assign v_G2_6447_out0 = v_RD_3283_out0 && v_RM_5974_out0;
assign v_CARRY_2784_out0 = v_G2_6447_out0;
assign v_S_4771_out0 = v_G1_4202_out0;
assign v_S_795_out0 = v_S_4771_out0;
assign v_G1_2147_out0 = v_CARRY_2784_out0 || v_CARRY_2783_out0;
assign v_COUT_531_out0 = v_G1_2147_out0;
assign v__3465_out0 = { v__1257_out0,v_S_795_out0 };
assign v_CIN_5030_out0 = v_COUT_531_out0;
assign v_RD_3281_out0 = v_CIN_5030_out0;
assign v_G1_4200_out0 = ((v_RD_3281_out0 && !v_RM_5972_out0) || (!v_RD_3281_out0) && v_RM_5972_out0);
assign v_G2_6445_out0 = v_RD_3281_out0 && v_RM_5972_out0;
assign v_CARRY_2782_out0 = v_G2_6445_out0;
assign v_S_4769_out0 = v_G1_4200_out0;
assign v_S_794_out0 = v_S_4769_out0;
assign v_G1_2146_out0 = v_CARRY_2782_out0 || v_CARRY_2781_out0;
assign v_COUT_530_out0 = v_G1_2146_out0;
assign v__6675_out0 = { v__3465_out0,v_S_794_out0 };
assign v_CIN_5037_out0 = v_COUT_530_out0;
assign v_RD_3296_out0 = v_CIN_5037_out0;
assign v_G1_4215_out0 = ((v_RD_3296_out0 && !v_RM_5987_out0) || (!v_RD_3296_out0) && v_RM_5987_out0);
assign v_G2_6460_out0 = v_RD_3296_out0 && v_RM_5987_out0;
assign v_CARRY_2797_out0 = v_G2_6460_out0;
assign v_S_4784_out0 = v_G1_4215_out0;
assign v_S_801_out0 = v_S_4784_out0;
assign v_G1_2153_out0 = v_CARRY_2797_out0 || v_CARRY_2796_out0;
assign v_COUT_537_out0 = v_G1_2153_out0;
assign v__1623_out0 = { v__6675_out0,v_S_801_out0 };
assign v_CIN_5038_out0 = v_COUT_537_out0;
assign v_RD_3298_out0 = v_CIN_5038_out0;
assign v_G1_4217_out0 = ((v_RD_3298_out0 && !v_RM_5989_out0) || (!v_RD_3298_out0) && v_RM_5989_out0);
assign v_G2_6462_out0 = v_RD_3298_out0 && v_RM_5989_out0;
assign v_CARRY_2799_out0 = v_G2_6462_out0;
assign v_S_4786_out0 = v_G1_4217_out0;
assign v_S_802_out0 = v_S_4786_out0;
assign v_G1_2154_out0 = v_CARRY_2799_out0 || v_CARRY_2798_out0;
assign v_COUT_538_out0 = v_G1_2154_out0;
assign v__3520_out0 = { v__1623_out0,v_S_802_out0 };
assign v_CIN_5040_out0 = v_COUT_538_out0;
assign v_RD_3302_out0 = v_CIN_5040_out0;
assign v_G1_4221_out0 = ((v_RD_3302_out0 && !v_RM_5993_out0) || (!v_RD_3302_out0) && v_RM_5993_out0);
assign v_G2_6466_out0 = v_RD_3302_out0 && v_RM_5993_out0;
assign v_CARRY_2803_out0 = v_G2_6466_out0;
assign v_S_4790_out0 = v_G1_4221_out0;
assign v_S_804_out0 = v_S_4790_out0;
assign v_G1_2156_out0 = v_CARRY_2803_out0 || v_CARRY_2802_out0;
assign v_COUT_540_out0 = v_G1_2156_out0;
assign v__2331_out0 = { v__3520_out0,v_S_804_out0 };
assign v_CIN_5033_out0 = v_COUT_540_out0;
assign v_RD_3288_out0 = v_CIN_5033_out0;
assign v_G1_4207_out0 = ((v_RD_3288_out0 && !v_RM_5979_out0) || (!v_RD_3288_out0) && v_RM_5979_out0);
assign v_G2_6452_out0 = v_RD_3288_out0 && v_RM_5979_out0;
assign v_CARRY_2789_out0 = v_G2_6452_out0;
assign v_S_4776_out0 = v_G1_4207_out0;
assign v_S_797_out0 = v_S_4776_out0;
assign v_G1_2149_out0 = v_CARRY_2789_out0 || v_CARRY_2788_out0;
assign v_COUT_533_out0 = v_G1_2149_out0;
assign v__3413_out0 = { v__2331_out0,v_S_797_out0 };
assign v_CIN_5034_out0 = v_COUT_533_out0;
assign v_RD_3290_out0 = v_CIN_5034_out0;
assign v_G1_4209_out0 = ((v_RD_3290_out0 && !v_RM_5981_out0) || (!v_RD_3290_out0) && v_RM_5981_out0);
assign v_G2_6454_out0 = v_RD_3290_out0 && v_RM_5981_out0;
assign v_CARRY_2791_out0 = v_G2_6454_out0;
assign v_S_4778_out0 = v_G1_4209_out0;
assign v_S_798_out0 = v_S_4778_out0;
assign v_G1_2150_out0 = v_CARRY_2791_out0 || v_CARRY_2790_out0;
assign v_COUT_534_out0 = v_G1_2150_out0;
assign v__2857_out0 = { v__3413_out0,v_S_798_out0 };
assign v_CIN_5039_out0 = v_COUT_534_out0;
assign v_RD_3300_out0 = v_CIN_5039_out0;
assign v_G1_4219_out0 = ((v_RD_3300_out0 && !v_RM_5991_out0) || (!v_RD_3300_out0) && v_RM_5991_out0);
assign v_G2_6464_out0 = v_RD_3300_out0 && v_RM_5991_out0;
assign v_CARRY_2801_out0 = v_G2_6464_out0;
assign v_S_4788_out0 = v_G1_4219_out0;
assign v_S_803_out0 = v_S_4788_out0;
assign v_G1_2155_out0 = v_CARRY_2801_out0 || v_CARRY_2800_out0;
assign v_COUT_539_out0 = v_G1_2155_out0;
assign v__1001_out0 = { v__2857_out0,v_S_803_out0 };
assign v_CIN_5027_out0 = v_COUT_539_out0;
assign v_RD_3275_out0 = v_CIN_5027_out0;
assign v_G1_4194_out0 = ((v_RD_3275_out0 && !v_RM_5966_out0) || (!v_RD_3275_out0) && v_RM_5966_out0);
assign v_G2_6439_out0 = v_RD_3275_out0 && v_RM_5966_out0;
assign v_CARRY_2776_out0 = v_G2_6439_out0;
assign v_S_4763_out0 = v_G1_4194_out0;
assign v_S_791_out0 = v_S_4763_out0;
assign v_G1_2143_out0 = v_CARRY_2776_out0 || v_CARRY_2775_out0;
assign v_COUT_527_out0 = v_G1_2143_out0;
assign v__1377_out0 = { v__1001_out0,v_S_791_out0 };
assign v_CIN_5032_out0 = v_COUT_527_out0;
assign v_RD_3285_out0 = v_CIN_5032_out0;
assign v_G1_4204_out0 = ((v_RD_3285_out0 && !v_RM_5976_out0) || (!v_RD_3285_out0) && v_RM_5976_out0);
assign v_G2_6449_out0 = v_RD_3285_out0 && v_RM_5976_out0;
assign v_CARRY_2786_out0 = v_G2_6449_out0;
assign v_S_4773_out0 = v_G1_4204_out0;
assign v_S_796_out0 = v_S_4773_out0;
assign v_G1_2148_out0 = v_CARRY_2786_out0 || v_CARRY_2785_out0;
assign v_COUT_532_out0 = v_G1_2148_out0;
assign v__904_out0 = { v__1377_out0,v_S_796_out0 };
assign v_CIN_5028_out0 = v_COUT_532_out0;
assign v_RD_3277_out0 = v_CIN_5028_out0;
assign v_G1_4196_out0 = ((v_RD_3277_out0 && !v_RM_5968_out0) || (!v_RD_3277_out0) && v_RM_5968_out0);
assign v_G2_6441_out0 = v_RD_3277_out0 && v_RM_5968_out0;
assign v_CARRY_2778_out0 = v_G2_6441_out0;
assign v_S_4765_out0 = v_G1_4196_out0;
assign v_S_792_out0 = v_S_4765_out0;
assign v_G1_2144_out0 = v_CARRY_2778_out0 || v_CARRY_2777_out0;
assign v_COUT_528_out0 = v_G1_2144_out0;
assign v__2233_out0 = { v__904_out0,v_S_792_out0 };
assign v_RM_1826_out0 = v_COUT_528_out0;
assign v_RM_5969_out0 = v_RM_1826_out0;
assign v_G1_4197_out0 = ((v_RD_3278_out0 && !v_RM_5969_out0) || (!v_RD_3278_out0) && v_RM_5969_out0);
assign v_G2_6442_out0 = v_RD_3278_out0 && v_RM_5969_out0;
assign v_CARRY_2779_out0 = v_G2_6442_out0;
assign v_S_4766_out0 = v_G1_4197_out0;
assign v_RM_5970_out0 = v_S_4766_out0;
assign v_G1_4198_out0 = ((v_RD_3279_out0 && !v_RM_5970_out0) || (!v_RD_3279_out0) && v_RM_5970_out0);
assign v_G2_6443_out0 = v_RD_3279_out0 && v_RM_5970_out0;
assign v_CARRY_2780_out0 = v_G2_6443_out0;
assign v_S_4767_out0 = v_G1_4198_out0;
assign v_S_793_out0 = v_S_4767_out0;
assign v_G1_2145_out0 = v_CARRY_2780_out0 || v_CARRY_2779_out0;
assign v_COUT_529_out0 = v_G1_2145_out0;
assign v__5256_out0 = { v__2233_out0,v_S_793_out0 };
assign v__5399_out0 = { v__5256_out0,v_COUT_529_out0 };
assign v_COUT_5384_out0 = v__5399_out0;
assign v_CIN_1158_out0 = v_COUT_5384_out0;
assign v__240_out0 = v_CIN_1158_out0[8:8];
assign v__878_out0 = v_CIN_1158_out0[6:6];
assign v__1061_out0 = v_CIN_1158_out0[3:3];
assign v__1080_out0 = v_CIN_1158_out0[15:15];
assign v__1231_out0 = v_CIN_1158_out0[0:0];
assign v__1499_out0 = v_CIN_1158_out0[9:9];
assign v__1515_out0 = v_CIN_1158_out0[2:2];
assign v__1541_out0 = v_CIN_1158_out0[7:7];
assign v__1874_out0 = v_CIN_1158_out0[1:1];
assign v__1892_out0 = v_CIN_1158_out0[10:10];
assign v__3351_out0 = v_CIN_1158_out0[11:11];
assign v__3767_out0 = v_CIN_1158_out0[12:12];
assign v__4293_out0 = v_CIN_1158_out0[13:13];
assign v__4326_out0 = v_CIN_1158_out0[14:14];
assign v__5287_out0 = v_CIN_1158_out0[5:5];
assign v__6635_out0 = v_CIN_1158_out0[4:4];
assign v_RM_1794_out0 = v__3767_out0;
assign v_RM_1795_out0 = v__4326_out0;
assign v_RM_1797_out0 = v__5287_out0;
assign v_RM_1798_out0 = v__6635_out0;
assign v_RM_1799_out0 = v__4293_out0;
assign v_RM_1800_out0 = v__1499_out0;
assign v_RM_1801_out0 = v__1892_out0;
assign v_RM_1802_out0 = v__1874_out0;
assign v_RM_1803_out0 = v__1061_out0;
assign v_RM_1804_out0 = v__878_out0;
assign v_RM_1805_out0 = v__1541_out0;
assign v_RM_1806_out0 = v__3351_out0;
assign v_RM_1807_out0 = v__240_out0;
assign v_RM_1808_out0 = v__1515_out0;
assign v_CIN_4999_out0 = v__1080_out0;
assign v_RM_5915_out0 = v__1231_out0;
assign v_RD_3217_out0 = v_CIN_4999_out0;
assign v_G1_4143_out0 = ((v_RD_3224_out0 && !v_RM_5915_out0) || (!v_RD_3224_out0) && v_RM_5915_out0);
assign v_RM_5903_out0 = v_RM_1794_out0;
assign v_RM_5905_out0 = v_RM_1795_out0;
assign v_RM_5909_out0 = v_RM_1797_out0;
assign v_RM_5911_out0 = v_RM_1798_out0;
assign v_RM_5913_out0 = v_RM_1799_out0;
assign v_RM_5916_out0 = v_RM_1800_out0;
assign v_RM_5918_out0 = v_RM_1801_out0;
assign v_RM_5920_out0 = v_RM_1802_out0;
assign v_RM_5922_out0 = v_RM_1803_out0;
assign v_RM_5924_out0 = v_RM_1804_out0;
assign v_RM_5926_out0 = v_RM_1805_out0;
assign v_RM_5928_out0 = v_RM_1806_out0;
assign v_RM_5930_out0 = v_RM_1807_out0;
assign v_RM_5932_out0 = v_RM_1808_out0;
assign v_G2_6388_out0 = v_RD_3224_out0 && v_RM_5915_out0;
assign v_CARRY_2725_out0 = v_G2_6388_out0;
assign v_G1_4131_out0 = ((v_RD_3212_out0 && !v_RM_5903_out0) || (!v_RD_3212_out0) && v_RM_5903_out0);
assign v_G1_4133_out0 = ((v_RD_3214_out0 && !v_RM_5905_out0) || (!v_RD_3214_out0) && v_RM_5905_out0);
assign v_G1_4137_out0 = ((v_RD_3218_out0 && !v_RM_5909_out0) || (!v_RD_3218_out0) && v_RM_5909_out0);
assign v_G1_4139_out0 = ((v_RD_3220_out0 && !v_RM_5911_out0) || (!v_RD_3220_out0) && v_RM_5911_out0);
assign v_G1_4141_out0 = ((v_RD_3222_out0 && !v_RM_5913_out0) || (!v_RD_3222_out0) && v_RM_5913_out0);
assign v_G1_4144_out0 = ((v_RD_3225_out0 && !v_RM_5916_out0) || (!v_RD_3225_out0) && v_RM_5916_out0);
assign v_G1_4146_out0 = ((v_RD_3227_out0 && !v_RM_5918_out0) || (!v_RD_3227_out0) && v_RM_5918_out0);
assign v_G1_4148_out0 = ((v_RD_3229_out0 && !v_RM_5920_out0) || (!v_RD_3229_out0) && v_RM_5920_out0);
assign v_G1_4150_out0 = ((v_RD_3231_out0 && !v_RM_5922_out0) || (!v_RD_3231_out0) && v_RM_5922_out0);
assign v_G1_4152_out0 = ((v_RD_3233_out0 && !v_RM_5924_out0) || (!v_RD_3233_out0) && v_RM_5924_out0);
assign v_G1_4154_out0 = ((v_RD_3235_out0 && !v_RM_5926_out0) || (!v_RD_3235_out0) && v_RM_5926_out0);
assign v_G1_4156_out0 = ((v_RD_3237_out0 && !v_RM_5928_out0) || (!v_RD_3237_out0) && v_RM_5928_out0);
assign v_G1_4158_out0 = ((v_RD_3239_out0 && !v_RM_5930_out0) || (!v_RD_3239_out0) && v_RM_5930_out0);
assign v_G1_4160_out0 = ((v_RD_3241_out0 && !v_RM_5932_out0) || (!v_RD_3241_out0) && v_RM_5932_out0);
assign v_S_4712_out0 = v_G1_4143_out0;
assign v_G2_6376_out0 = v_RD_3212_out0 && v_RM_5903_out0;
assign v_G2_6378_out0 = v_RD_3214_out0 && v_RM_5905_out0;
assign v_G2_6382_out0 = v_RD_3218_out0 && v_RM_5909_out0;
assign v_G2_6384_out0 = v_RD_3220_out0 && v_RM_5911_out0;
assign v_G2_6386_out0 = v_RD_3222_out0 && v_RM_5913_out0;
assign v_G2_6389_out0 = v_RD_3225_out0 && v_RM_5916_out0;
assign v_G2_6391_out0 = v_RD_3227_out0 && v_RM_5918_out0;
assign v_G2_6393_out0 = v_RD_3229_out0 && v_RM_5920_out0;
assign v_G2_6395_out0 = v_RD_3231_out0 && v_RM_5922_out0;
assign v_G2_6397_out0 = v_RD_3233_out0 && v_RM_5924_out0;
assign v_G2_6399_out0 = v_RD_3235_out0 && v_RM_5926_out0;
assign v_G2_6401_out0 = v_RD_3237_out0 && v_RM_5928_out0;
assign v_G2_6403_out0 = v_RD_3239_out0 && v_RM_5930_out0;
assign v_G2_6405_out0 = v_RD_3241_out0 && v_RM_5932_out0;
assign v_S_2289_out0 = v_S_4712_out0;
assign v_CARRY_2713_out0 = v_G2_6376_out0;
assign v_CARRY_2715_out0 = v_G2_6378_out0;
assign v_CARRY_2719_out0 = v_G2_6382_out0;
assign v_CARRY_2721_out0 = v_G2_6384_out0;
assign v_CARRY_2723_out0 = v_G2_6386_out0;
assign v_CARRY_2726_out0 = v_G2_6389_out0;
assign v_CARRY_2728_out0 = v_G2_6391_out0;
assign v_CARRY_2730_out0 = v_G2_6393_out0;
assign v_CARRY_2732_out0 = v_G2_6395_out0;
assign v_CARRY_2734_out0 = v_G2_6397_out0;
assign v_CARRY_2736_out0 = v_G2_6399_out0;
assign v_CARRY_2738_out0 = v_G2_6401_out0;
assign v_CARRY_2740_out0 = v_G2_6403_out0;
assign v_CARRY_2742_out0 = v_G2_6405_out0;
assign v_S_4700_out0 = v_G1_4131_out0;
assign v_S_4702_out0 = v_G1_4133_out0;
assign v_S_4706_out0 = v_G1_4137_out0;
assign v_S_4708_out0 = v_G1_4139_out0;
assign v_S_4710_out0 = v_G1_4141_out0;
assign v_S_4713_out0 = v_G1_4144_out0;
assign v_S_4715_out0 = v_G1_4146_out0;
assign v_S_4717_out0 = v_G1_4148_out0;
assign v_S_4719_out0 = v_G1_4150_out0;
assign v_S_4721_out0 = v_G1_4152_out0;
assign v_S_4723_out0 = v_G1_4154_out0;
assign v_S_4725_out0 = v_G1_4156_out0;
assign v_S_4727_out0 = v_G1_4158_out0;
assign v_S_4729_out0 = v_G1_4160_out0;
assign v_CIN_5005_out0 = v_CARRY_2725_out0;
assign v__308_out0 = { v__330_out0,v_S_2289_out0 };
assign v_RD_3230_out0 = v_CIN_5005_out0;
assign v_RM_5904_out0 = v_S_4700_out0;
assign v_RM_5906_out0 = v_S_4702_out0;
assign v_RM_5910_out0 = v_S_4706_out0;
assign v_RM_5912_out0 = v_S_4708_out0;
assign v_RM_5914_out0 = v_S_4710_out0;
assign v_RM_5917_out0 = v_S_4713_out0;
assign v_RM_5919_out0 = v_S_4715_out0;
assign v_RM_5921_out0 = v_S_4717_out0;
assign v_RM_5923_out0 = v_S_4719_out0;
assign v_RM_5925_out0 = v_S_4721_out0;
assign v_RM_5927_out0 = v_S_4723_out0;
assign v_RM_5929_out0 = v_S_4725_out0;
assign v_RM_5931_out0 = v_S_4727_out0;
assign v_RM_5933_out0 = v_S_4729_out0;
assign v_G1_4149_out0 = ((v_RD_3230_out0 && !v_RM_5921_out0) || (!v_RD_3230_out0) && v_RM_5921_out0);
assign v_G2_6394_out0 = v_RD_3230_out0 && v_RM_5921_out0;
assign v_CARRY_2731_out0 = v_G2_6394_out0;
assign v_S_4718_out0 = v_G1_4149_out0;
assign v_S_769_out0 = v_S_4718_out0;
assign v_G1_2121_out0 = v_CARRY_2731_out0 || v_CARRY_2730_out0;
assign v_COUT_505_out0 = v_G1_2121_out0;
assign v_CIN_5011_out0 = v_COUT_505_out0;
assign v_RD_3242_out0 = v_CIN_5011_out0;
assign v_G1_4161_out0 = ((v_RD_3242_out0 && !v_RM_5933_out0) || (!v_RD_3242_out0) && v_RM_5933_out0);
assign v_G2_6406_out0 = v_RD_3242_out0 && v_RM_5933_out0;
assign v_CARRY_2743_out0 = v_G2_6406_out0;
assign v_S_4730_out0 = v_G1_4161_out0;
assign v_S_775_out0 = v_S_4730_out0;
assign v_G1_2127_out0 = v_CARRY_2743_out0 || v_CARRY_2742_out0;
assign v_COUT_511_out0 = v_G1_2127_out0;
assign v__2346_out0 = { v_S_769_out0,v_S_775_out0 };
assign v_CIN_5006_out0 = v_COUT_511_out0;
assign v_RD_3232_out0 = v_CIN_5006_out0;
assign v_G1_4151_out0 = ((v_RD_3232_out0 && !v_RM_5923_out0) || (!v_RD_3232_out0) && v_RM_5923_out0);
assign v_G2_6396_out0 = v_RD_3232_out0 && v_RM_5923_out0;
assign v_CARRY_2733_out0 = v_G2_6396_out0;
assign v_S_4720_out0 = v_G1_4151_out0;
assign v_S_770_out0 = v_S_4720_out0;
assign v_G1_2122_out0 = v_CARRY_2733_out0 || v_CARRY_2732_out0;
assign v_COUT_506_out0 = v_G1_2122_out0;
assign v__1255_out0 = { v__2346_out0,v_S_770_out0 };
assign v_CIN_5001_out0 = v_COUT_506_out0;
assign v_RD_3221_out0 = v_CIN_5001_out0;
assign v_G1_4140_out0 = ((v_RD_3221_out0 && !v_RM_5912_out0) || (!v_RD_3221_out0) && v_RM_5912_out0);
assign v_G2_6385_out0 = v_RD_3221_out0 && v_RM_5912_out0;
assign v_CARRY_2722_out0 = v_G2_6385_out0;
assign v_S_4709_out0 = v_G1_4140_out0;
assign v_S_765_out0 = v_S_4709_out0;
assign v_G1_2117_out0 = v_CARRY_2722_out0 || v_CARRY_2721_out0;
assign v_COUT_501_out0 = v_G1_2117_out0;
assign v__3463_out0 = { v__1255_out0,v_S_765_out0 };
assign v_CIN_5000_out0 = v_COUT_501_out0;
assign v_RD_3219_out0 = v_CIN_5000_out0;
assign v_G1_4138_out0 = ((v_RD_3219_out0 && !v_RM_5910_out0) || (!v_RD_3219_out0) && v_RM_5910_out0);
assign v_G2_6383_out0 = v_RD_3219_out0 && v_RM_5910_out0;
assign v_CARRY_2720_out0 = v_G2_6383_out0;
assign v_S_4707_out0 = v_G1_4138_out0;
assign v_S_764_out0 = v_S_4707_out0;
assign v_G1_2116_out0 = v_CARRY_2720_out0 || v_CARRY_2719_out0;
assign v_COUT_500_out0 = v_G1_2116_out0;
assign v__6673_out0 = { v__3463_out0,v_S_764_out0 };
assign v_CIN_5007_out0 = v_COUT_500_out0;
assign v_RD_3234_out0 = v_CIN_5007_out0;
assign v_G1_4153_out0 = ((v_RD_3234_out0 && !v_RM_5925_out0) || (!v_RD_3234_out0) && v_RM_5925_out0);
assign v_G2_6398_out0 = v_RD_3234_out0 && v_RM_5925_out0;
assign v_CARRY_2735_out0 = v_G2_6398_out0;
assign v_S_4722_out0 = v_G1_4153_out0;
assign v_S_771_out0 = v_S_4722_out0;
assign v_G1_2123_out0 = v_CARRY_2735_out0 || v_CARRY_2734_out0;
assign v_COUT_507_out0 = v_G1_2123_out0;
assign v__1621_out0 = { v__6673_out0,v_S_771_out0 };
assign v_CIN_5008_out0 = v_COUT_507_out0;
assign v_RD_3236_out0 = v_CIN_5008_out0;
assign v_G1_4155_out0 = ((v_RD_3236_out0 && !v_RM_5927_out0) || (!v_RD_3236_out0) && v_RM_5927_out0);
assign v_G2_6400_out0 = v_RD_3236_out0 && v_RM_5927_out0;
assign v_CARRY_2737_out0 = v_G2_6400_out0;
assign v_S_4724_out0 = v_G1_4155_out0;
assign v_S_772_out0 = v_S_4724_out0;
assign v_G1_2124_out0 = v_CARRY_2737_out0 || v_CARRY_2736_out0;
assign v_COUT_508_out0 = v_G1_2124_out0;
assign v__3518_out0 = { v__1621_out0,v_S_772_out0 };
assign v_CIN_5010_out0 = v_COUT_508_out0;
assign v_RD_3240_out0 = v_CIN_5010_out0;
assign v_G1_4159_out0 = ((v_RD_3240_out0 && !v_RM_5931_out0) || (!v_RD_3240_out0) && v_RM_5931_out0);
assign v_G2_6404_out0 = v_RD_3240_out0 && v_RM_5931_out0;
assign v_CARRY_2741_out0 = v_G2_6404_out0;
assign v_S_4728_out0 = v_G1_4159_out0;
assign v_S_774_out0 = v_S_4728_out0;
assign v_G1_2126_out0 = v_CARRY_2741_out0 || v_CARRY_2740_out0;
assign v_COUT_510_out0 = v_G1_2126_out0;
assign v__2329_out0 = { v__3518_out0,v_S_774_out0 };
assign v_CIN_5003_out0 = v_COUT_510_out0;
assign v_RD_3226_out0 = v_CIN_5003_out0;
assign v_G1_4145_out0 = ((v_RD_3226_out0 && !v_RM_5917_out0) || (!v_RD_3226_out0) && v_RM_5917_out0);
assign v_G2_6390_out0 = v_RD_3226_out0 && v_RM_5917_out0;
assign v_CARRY_2727_out0 = v_G2_6390_out0;
assign v_S_4714_out0 = v_G1_4145_out0;
assign v_S_767_out0 = v_S_4714_out0;
assign v_G1_2119_out0 = v_CARRY_2727_out0 || v_CARRY_2726_out0;
assign v_COUT_503_out0 = v_G1_2119_out0;
assign v__3411_out0 = { v__2329_out0,v_S_767_out0 };
assign v_CIN_5004_out0 = v_COUT_503_out0;
assign v_RD_3228_out0 = v_CIN_5004_out0;
assign v_G1_4147_out0 = ((v_RD_3228_out0 && !v_RM_5919_out0) || (!v_RD_3228_out0) && v_RM_5919_out0);
assign v_G2_6392_out0 = v_RD_3228_out0 && v_RM_5919_out0;
assign v_CARRY_2729_out0 = v_G2_6392_out0;
assign v_S_4716_out0 = v_G1_4147_out0;
assign v_S_768_out0 = v_S_4716_out0;
assign v_G1_2120_out0 = v_CARRY_2729_out0 || v_CARRY_2728_out0;
assign v_COUT_504_out0 = v_G1_2120_out0;
assign v__2855_out0 = { v__3411_out0,v_S_768_out0 };
assign v_CIN_5009_out0 = v_COUT_504_out0;
assign v_RD_3238_out0 = v_CIN_5009_out0;
assign v_G1_4157_out0 = ((v_RD_3238_out0 && !v_RM_5929_out0) || (!v_RD_3238_out0) && v_RM_5929_out0);
assign v_G2_6402_out0 = v_RD_3238_out0 && v_RM_5929_out0;
assign v_CARRY_2739_out0 = v_G2_6402_out0;
assign v_S_4726_out0 = v_G1_4157_out0;
assign v_S_773_out0 = v_S_4726_out0;
assign v_G1_2125_out0 = v_CARRY_2739_out0 || v_CARRY_2738_out0;
assign v_COUT_509_out0 = v_G1_2125_out0;
assign v__999_out0 = { v__2855_out0,v_S_773_out0 };
assign v_CIN_4997_out0 = v_COUT_509_out0;
assign v_RD_3213_out0 = v_CIN_4997_out0;
assign v_G1_4132_out0 = ((v_RD_3213_out0 && !v_RM_5904_out0) || (!v_RD_3213_out0) && v_RM_5904_out0);
assign v_G2_6377_out0 = v_RD_3213_out0 && v_RM_5904_out0;
assign v_CARRY_2714_out0 = v_G2_6377_out0;
assign v_S_4701_out0 = v_G1_4132_out0;
assign v_S_761_out0 = v_S_4701_out0;
assign v_G1_2113_out0 = v_CARRY_2714_out0 || v_CARRY_2713_out0;
assign v_COUT_497_out0 = v_G1_2113_out0;
assign v__1375_out0 = { v__999_out0,v_S_761_out0 };
assign v_CIN_5002_out0 = v_COUT_497_out0;
assign v_RD_3223_out0 = v_CIN_5002_out0;
assign v_G1_4142_out0 = ((v_RD_3223_out0 && !v_RM_5914_out0) || (!v_RD_3223_out0) && v_RM_5914_out0);
assign v_G2_6387_out0 = v_RD_3223_out0 && v_RM_5914_out0;
assign v_CARRY_2724_out0 = v_G2_6387_out0;
assign v_S_4711_out0 = v_G1_4142_out0;
assign v_S_766_out0 = v_S_4711_out0;
assign v_G1_2118_out0 = v_CARRY_2724_out0 || v_CARRY_2723_out0;
assign v_COUT_502_out0 = v_G1_2118_out0;
assign v__902_out0 = { v__1375_out0,v_S_766_out0 };
assign v_CIN_4998_out0 = v_COUT_502_out0;
assign v_RD_3215_out0 = v_CIN_4998_out0;
assign v_G1_4134_out0 = ((v_RD_3215_out0 && !v_RM_5906_out0) || (!v_RD_3215_out0) && v_RM_5906_out0);
assign v_G2_6379_out0 = v_RD_3215_out0 && v_RM_5906_out0;
assign v_CARRY_2716_out0 = v_G2_6379_out0;
assign v_S_4703_out0 = v_G1_4134_out0;
assign v_S_762_out0 = v_S_4703_out0;
assign v_G1_2114_out0 = v_CARRY_2716_out0 || v_CARRY_2715_out0;
assign v_COUT_498_out0 = v_G1_2114_out0;
assign v__2231_out0 = { v__902_out0,v_S_762_out0 };
assign v_RM_1796_out0 = v_COUT_498_out0;
assign v_RM_5907_out0 = v_RM_1796_out0;
assign v_G1_4135_out0 = ((v_RD_3216_out0 && !v_RM_5907_out0) || (!v_RD_3216_out0) && v_RM_5907_out0);
assign v_G2_6380_out0 = v_RD_3216_out0 && v_RM_5907_out0;
assign v_CARRY_2717_out0 = v_G2_6380_out0;
assign v_S_4704_out0 = v_G1_4135_out0;
assign v_RM_5908_out0 = v_S_4704_out0;
assign v_G1_4136_out0 = ((v_RD_3217_out0 && !v_RM_5908_out0) || (!v_RD_3217_out0) && v_RM_5908_out0);
assign v_G2_6381_out0 = v_RD_3217_out0 && v_RM_5908_out0;
assign v_CARRY_2718_out0 = v_G2_6381_out0;
assign v_S_4705_out0 = v_G1_4136_out0;
assign v_S_763_out0 = v_S_4705_out0;
assign v_G1_2115_out0 = v_CARRY_2718_out0 || v_CARRY_2717_out0;
assign v_COUT_499_out0 = v_G1_2115_out0;
assign v__5254_out0 = { v__2231_out0,v_S_763_out0 };
assign v__5397_out0 = { v__5254_out0,v_COUT_499_out0 };
assign v_COUT_5382_out0 = v__5397_out0;
assign v_CIN_1156_out0 = v_COUT_5382_out0;
assign v__238_out0 = v_CIN_1156_out0[8:8];
assign v__876_out0 = v_CIN_1156_out0[6:6];
assign v__1059_out0 = v_CIN_1156_out0[3:3];
assign v__1078_out0 = v_CIN_1156_out0[15:15];
assign v__1229_out0 = v_CIN_1156_out0[0:0];
assign v__1497_out0 = v_CIN_1156_out0[9:9];
assign v__1513_out0 = v_CIN_1156_out0[2:2];
assign v__1539_out0 = v_CIN_1156_out0[7:7];
assign v__1872_out0 = v_CIN_1156_out0[1:1];
assign v__1890_out0 = v_CIN_1156_out0[10:10];
assign v__3349_out0 = v_CIN_1156_out0[11:11];
assign v__3765_out0 = v_CIN_1156_out0[12:12];
assign v__4291_out0 = v_CIN_1156_out0[13:13];
assign v__4324_out0 = v_CIN_1156_out0[14:14];
assign v__5285_out0 = v_CIN_1156_out0[5:5];
assign v__6633_out0 = v_CIN_1156_out0[4:4];
assign v_RM_1764_out0 = v__3765_out0;
assign v_RM_1765_out0 = v__4324_out0;
assign v_RM_1767_out0 = v__5285_out0;
assign v_RM_1768_out0 = v__6633_out0;
assign v_RM_1769_out0 = v__4291_out0;
assign v_RM_1770_out0 = v__1497_out0;
assign v_RM_1771_out0 = v__1890_out0;
assign v_RM_1772_out0 = v__1872_out0;
assign v_RM_1773_out0 = v__1059_out0;
assign v_RM_1774_out0 = v__876_out0;
assign v_RM_1775_out0 = v__1539_out0;
assign v_RM_1776_out0 = v__3349_out0;
assign v_RM_1777_out0 = v__238_out0;
assign v_RM_1778_out0 = v__1513_out0;
assign v_CIN_4969_out0 = v__1078_out0;
assign v_RM_5853_out0 = v__1229_out0;
assign v_RD_3155_out0 = v_CIN_4969_out0;
assign v_G1_4081_out0 = ((v_RD_3162_out0 && !v_RM_5853_out0) || (!v_RD_3162_out0) && v_RM_5853_out0);
assign v_RM_5841_out0 = v_RM_1764_out0;
assign v_RM_5843_out0 = v_RM_1765_out0;
assign v_RM_5847_out0 = v_RM_1767_out0;
assign v_RM_5849_out0 = v_RM_1768_out0;
assign v_RM_5851_out0 = v_RM_1769_out0;
assign v_RM_5854_out0 = v_RM_1770_out0;
assign v_RM_5856_out0 = v_RM_1771_out0;
assign v_RM_5858_out0 = v_RM_1772_out0;
assign v_RM_5860_out0 = v_RM_1773_out0;
assign v_RM_5862_out0 = v_RM_1774_out0;
assign v_RM_5864_out0 = v_RM_1775_out0;
assign v_RM_5866_out0 = v_RM_1776_out0;
assign v_RM_5868_out0 = v_RM_1777_out0;
assign v_RM_5870_out0 = v_RM_1778_out0;
assign v_G2_6326_out0 = v_RD_3162_out0 && v_RM_5853_out0;
assign v_CARRY_2663_out0 = v_G2_6326_out0;
assign v_G1_4069_out0 = ((v_RD_3150_out0 && !v_RM_5841_out0) || (!v_RD_3150_out0) && v_RM_5841_out0);
assign v_G1_4071_out0 = ((v_RD_3152_out0 && !v_RM_5843_out0) || (!v_RD_3152_out0) && v_RM_5843_out0);
assign v_G1_4075_out0 = ((v_RD_3156_out0 && !v_RM_5847_out0) || (!v_RD_3156_out0) && v_RM_5847_out0);
assign v_G1_4077_out0 = ((v_RD_3158_out0 && !v_RM_5849_out0) || (!v_RD_3158_out0) && v_RM_5849_out0);
assign v_G1_4079_out0 = ((v_RD_3160_out0 && !v_RM_5851_out0) || (!v_RD_3160_out0) && v_RM_5851_out0);
assign v_G1_4082_out0 = ((v_RD_3163_out0 && !v_RM_5854_out0) || (!v_RD_3163_out0) && v_RM_5854_out0);
assign v_G1_4084_out0 = ((v_RD_3165_out0 && !v_RM_5856_out0) || (!v_RD_3165_out0) && v_RM_5856_out0);
assign v_G1_4086_out0 = ((v_RD_3167_out0 && !v_RM_5858_out0) || (!v_RD_3167_out0) && v_RM_5858_out0);
assign v_G1_4088_out0 = ((v_RD_3169_out0 && !v_RM_5860_out0) || (!v_RD_3169_out0) && v_RM_5860_out0);
assign v_G1_4090_out0 = ((v_RD_3171_out0 && !v_RM_5862_out0) || (!v_RD_3171_out0) && v_RM_5862_out0);
assign v_G1_4092_out0 = ((v_RD_3173_out0 && !v_RM_5864_out0) || (!v_RD_3173_out0) && v_RM_5864_out0);
assign v_G1_4094_out0 = ((v_RD_3175_out0 && !v_RM_5866_out0) || (!v_RD_3175_out0) && v_RM_5866_out0);
assign v_G1_4096_out0 = ((v_RD_3177_out0 && !v_RM_5868_out0) || (!v_RD_3177_out0) && v_RM_5868_out0);
assign v_G1_4098_out0 = ((v_RD_3179_out0 && !v_RM_5870_out0) || (!v_RD_3179_out0) && v_RM_5870_out0);
assign v_S_4650_out0 = v_G1_4081_out0;
assign v_G2_6314_out0 = v_RD_3150_out0 && v_RM_5841_out0;
assign v_G2_6316_out0 = v_RD_3152_out0 && v_RM_5843_out0;
assign v_G2_6320_out0 = v_RD_3156_out0 && v_RM_5847_out0;
assign v_G2_6322_out0 = v_RD_3158_out0 && v_RM_5849_out0;
assign v_G2_6324_out0 = v_RD_3160_out0 && v_RM_5851_out0;
assign v_G2_6327_out0 = v_RD_3163_out0 && v_RM_5854_out0;
assign v_G2_6329_out0 = v_RD_3165_out0 && v_RM_5856_out0;
assign v_G2_6331_out0 = v_RD_3167_out0 && v_RM_5858_out0;
assign v_G2_6333_out0 = v_RD_3169_out0 && v_RM_5860_out0;
assign v_G2_6335_out0 = v_RD_3171_out0 && v_RM_5862_out0;
assign v_G2_6337_out0 = v_RD_3173_out0 && v_RM_5864_out0;
assign v_G2_6339_out0 = v_RD_3175_out0 && v_RM_5866_out0;
assign v_G2_6341_out0 = v_RD_3177_out0 && v_RM_5868_out0;
assign v_G2_6343_out0 = v_RD_3179_out0 && v_RM_5870_out0;
assign v_S_2287_out0 = v_S_4650_out0;
assign v_CARRY_2651_out0 = v_G2_6314_out0;
assign v_CARRY_2653_out0 = v_G2_6316_out0;
assign v_CARRY_2657_out0 = v_G2_6320_out0;
assign v_CARRY_2659_out0 = v_G2_6322_out0;
assign v_CARRY_2661_out0 = v_G2_6324_out0;
assign v_CARRY_2664_out0 = v_G2_6327_out0;
assign v_CARRY_2666_out0 = v_G2_6329_out0;
assign v_CARRY_2668_out0 = v_G2_6331_out0;
assign v_CARRY_2670_out0 = v_G2_6333_out0;
assign v_CARRY_2672_out0 = v_G2_6335_out0;
assign v_CARRY_2674_out0 = v_G2_6337_out0;
assign v_CARRY_2676_out0 = v_G2_6339_out0;
assign v_CARRY_2678_out0 = v_G2_6341_out0;
assign v_CARRY_2680_out0 = v_G2_6343_out0;
assign v_S_4638_out0 = v_G1_4069_out0;
assign v_S_4640_out0 = v_G1_4071_out0;
assign v_S_4644_out0 = v_G1_4075_out0;
assign v_S_4646_out0 = v_G1_4077_out0;
assign v_S_4648_out0 = v_G1_4079_out0;
assign v_S_4651_out0 = v_G1_4082_out0;
assign v_S_4653_out0 = v_G1_4084_out0;
assign v_S_4655_out0 = v_G1_4086_out0;
assign v_S_4657_out0 = v_G1_4088_out0;
assign v_S_4659_out0 = v_G1_4090_out0;
assign v_S_4661_out0 = v_G1_4092_out0;
assign v_S_4663_out0 = v_G1_4094_out0;
assign v_S_4665_out0 = v_G1_4096_out0;
assign v_S_4667_out0 = v_G1_4098_out0;
assign v_CIN_4975_out0 = v_CARRY_2663_out0;
assign v__24_out0 = { v__308_out0,v_S_2287_out0 };
assign v_RD_3168_out0 = v_CIN_4975_out0;
assign v_RM_5842_out0 = v_S_4638_out0;
assign v_RM_5844_out0 = v_S_4640_out0;
assign v_RM_5848_out0 = v_S_4644_out0;
assign v_RM_5850_out0 = v_S_4646_out0;
assign v_RM_5852_out0 = v_S_4648_out0;
assign v_RM_5855_out0 = v_S_4651_out0;
assign v_RM_5857_out0 = v_S_4653_out0;
assign v_RM_5859_out0 = v_S_4655_out0;
assign v_RM_5861_out0 = v_S_4657_out0;
assign v_RM_5863_out0 = v_S_4659_out0;
assign v_RM_5865_out0 = v_S_4661_out0;
assign v_RM_5867_out0 = v_S_4663_out0;
assign v_RM_5869_out0 = v_S_4665_out0;
assign v_RM_5871_out0 = v_S_4667_out0;
assign v_G1_4087_out0 = ((v_RD_3168_out0 && !v_RM_5859_out0) || (!v_RD_3168_out0) && v_RM_5859_out0);
assign v_G2_6332_out0 = v_RD_3168_out0 && v_RM_5859_out0;
assign v_CARRY_2669_out0 = v_G2_6332_out0;
assign v_S_4656_out0 = v_G1_4087_out0;
assign v_S_739_out0 = v_S_4656_out0;
assign v_G1_2091_out0 = v_CARRY_2669_out0 || v_CARRY_2668_out0;
assign v_COUT_475_out0 = v_G1_2091_out0;
assign v_CIN_4981_out0 = v_COUT_475_out0;
assign v_RD_3180_out0 = v_CIN_4981_out0;
assign v_G1_4099_out0 = ((v_RD_3180_out0 && !v_RM_5871_out0) || (!v_RD_3180_out0) && v_RM_5871_out0);
assign v_G2_6344_out0 = v_RD_3180_out0 && v_RM_5871_out0;
assign v_CARRY_2681_out0 = v_G2_6344_out0;
assign v_S_4668_out0 = v_G1_4099_out0;
assign v_S_745_out0 = v_S_4668_out0;
assign v_G1_2097_out0 = v_CARRY_2681_out0 || v_CARRY_2680_out0;
assign v_COUT_481_out0 = v_G1_2097_out0;
assign v__2344_out0 = { v_S_739_out0,v_S_745_out0 };
assign v_CIN_4976_out0 = v_COUT_481_out0;
assign v_RD_3170_out0 = v_CIN_4976_out0;
assign v_G1_4089_out0 = ((v_RD_3170_out0 && !v_RM_5861_out0) || (!v_RD_3170_out0) && v_RM_5861_out0);
assign v_G2_6334_out0 = v_RD_3170_out0 && v_RM_5861_out0;
assign v_CARRY_2671_out0 = v_G2_6334_out0;
assign v_S_4658_out0 = v_G1_4089_out0;
assign v_S_740_out0 = v_S_4658_out0;
assign v_G1_2092_out0 = v_CARRY_2671_out0 || v_CARRY_2670_out0;
assign v_COUT_476_out0 = v_G1_2092_out0;
assign v__1253_out0 = { v__2344_out0,v_S_740_out0 };
assign v_CIN_4971_out0 = v_COUT_476_out0;
assign v_RD_3159_out0 = v_CIN_4971_out0;
assign v_G1_4078_out0 = ((v_RD_3159_out0 && !v_RM_5850_out0) || (!v_RD_3159_out0) && v_RM_5850_out0);
assign v_G2_6323_out0 = v_RD_3159_out0 && v_RM_5850_out0;
assign v_CARRY_2660_out0 = v_G2_6323_out0;
assign v_S_4647_out0 = v_G1_4078_out0;
assign v_S_735_out0 = v_S_4647_out0;
assign v_G1_2087_out0 = v_CARRY_2660_out0 || v_CARRY_2659_out0;
assign v_COUT_471_out0 = v_G1_2087_out0;
assign v__3461_out0 = { v__1253_out0,v_S_735_out0 };
assign v_CIN_4970_out0 = v_COUT_471_out0;
assign v_RD_3157_out0 = v_CIN_4970_out0;
assign v_G1_4076_out0 = ((v_RD_3157_out0 && !v_RM_5848_out0) || (!v_RD_3157_out0) && v_RM_5848_out0);
assign v_G2_6321_out0 = v_RD_3157_out0 && v_RM_5848_out0;
assign v_CARRY_2658_out0 = v_G2_6321_out0;
assign v_S_4645_out0 = v_G1_4076_out0;
assign v_S_734_out0 = v_S_4645_out0;
assign v_G1_2086_out0 = v_CARRY_2658_out0 || v_CARRY_2657_out0;
assign v_COUT_470_out0 = v_G1_2086_out0;
assign v__6671_out0 = { v__3461_out0,v_S_734_out0 };
assign v_CIN_4977_out0 = v_COUT_470_out0;
assign v_RD_3172_out0 = v_CIN_4977_out0;
assign v_G1_4091_out0 = ((v_RD_3172_out0 && !v_RM_5863_out0) || (!v_RD_3172_out0) && v_RM_5863_out0);
assign v_G2_6336_out0 = v_RD_3172_out0 && v_RM_5863_out0;
assign v_CARRY_2673_out0 = v_G2_6336_out0;
assign v_S_4660_out0 = v_G1_4091_out0;
assign v_S_741_out0 = v_S_4660_out0;
assign v_G1_2093_out0 = v_CARRY_2673_out0 || v_CARRY_2672_out0;
assign v_COUT_477_out0 = v_G1_2093_out0;
assign v__1619_out0 = { v__6671_out0,v_S_741_out0 };
assign v_CIN_4978_out0 = v_COUT_477_out0;
assign v_RD_3174_out0 = v_CIN_4978_out0;
assign v_G1_4093_out0 = ((v_RD_3174_out0 && !v_RM_5865_out0) || (!v_RD_3174_out0) && v_RM_5865_out0);
assign v_G2_6338_out0 = v_RD_3174_out0 && v_RM_5865_out0;
assign v_CARRY_2675_out0 = v_G2_6338_out0;
assign v_S_4662_out0 = v_G1_4093_out0;
assign v_S_742_out0 = v_S_4662_out0;
assign v_G1_2094_out0 = v_CARRY_2675_out0 || v_CARRY_2674_out0;
assign v_COUT_478_out0 = v_G1_2094_out0;
assign v__3516_out0 = { v__1619_out0,v_S_742_out0 };
assign v_CIN_4980_out0 = v_COUT_478_out0;
assign v_RD_3178_out0 = v_CIN_4980_out0;
assign v_G1_4097_out0 = ((v_RD_3178_out0 && !v_RM_5869_out0) || (!v_RD_3178_out0) && v_RM_5869_out0);
assign v_G2_6342_out0 = v_RD_3178_out0 && v_RM_5869_out0;
assign v_CARRY_2679_out0 = v_G2_6342_out0;
assign v_S_4666_out0 = v_G1_4097_out0;
assign v_S_744_out0 = v_S_4666_out0;
assign v_G1_2096_out0 = v_CARRY_2679_out0 || v_CARRY_2678_out0;
assign v_COUT_480_out0 = v_G1_2096_out0;
assign v__2327_out0 = { v__3516_out0,v_S_744_out0 };
assign v_CIN_4973_out0 = v_COUT_480_out0;
assign v_RD_3164_out0 = v_CIN_4973_out0;
assign v_G1_4083_out0 = ((v_RD_3164_out0 && !v_RM_5855_out0) || (!v_RD_3164_out0) && v_RM_5855_out0);
assign v_G2_6328_out0 = v_RD_3164_out0 && v_RM_5855_out0;
assign v_CARRY_2665_out0 = v_G2_6328_out0;
assign v_S_4652_out0 = v_G1_4083_out0;
assign v_S_737_out0 = v_S_4652_out0;
assign v_G1_2089_out0 = v_CARRY_2665_out0 || v_CARRY_2664_out0;
assign v_COUT_473_out0 = v_G1_2089_out0;
assign v__3409_out0 = { v__2327_out0,v_S_737_out0 };
assign v_CIN_4974_out0 = v_COUT_473_out0;
assign v_RD_3166_out0 = v_CIN_4974_out0;
assign v_G1_4085_out0 = ((v_RD_3166_out0 && !v_RM_5857_out0) || (!v_RD_3166_out0) && v_RM_5857_out0);
assign v_G2_6330_out0 = v_RD_3166_out0 && v_RM_5857_out0;
assign v_CARRY_2667_out0 = v_G2_6330_out0;
assign v_S_4654_out0 = v_G1_4085_out0;
assign v_S_738_out0 = v_S_4654_out0;
assign v_G1_2090_out0 = v_CARRY_2667_out0 || v_CARRY_2666_out0;
assign v_COUT_474_out0 = v_G1_2090_out0;
assign v__2853_out0 = { v__3409_out0,v_S_738_out0 };
assign v_CIN_4979_out0 = v_COUT_474_out0;
assign v_RD_3176_out0 = v_CIN_4979_out0;
assign v_G1_4095_out0 = ((v_RD_3176_out0 && !v_RM_5867_out0) || (!v_RD_3176_out0) && v_RM_5867_out0);
assign v_G2_6340_out0 = v_RD_3176_out0 && v_RM_5867_out0;
assign v_CARRY_2677_out0 = v_G2_6340_out0;
assign v_S_4664_out0 = v_G1_4095_out0;
assign v_S_743_out0 = v_S_4664_out0;
assign v_G1_2095_out0 = v_CARRY_2677_out0 || v_CARRY_2676_out0;
assign v_COUT_479_out0 = v_G1_2095_out0;
assign v__997_out0 = { v__2853_out0,v_S_743_out0 };
assign v_CIN_4967_out0 = v_COUT_479_out0;
assign v_RD_3151_out0 = v_CIN_4967_out0;
assign v_G1_4070_out0 = ((v_RD_3151_out0 && !v_RM_5842_out0) || (!v_RD_3151_out0) && v_RM_5842_out0);
assign v_G2_6315_out0 = v_RD_3151_out0 && v_RM_5842_out0;
assign v_CARRY_2652_out0 = v_G2_6315_out0;
assign v_S_4639_out0 = v_G1_4070_out0;
assign v_S_731_out0 = v_S_4639_out0;
assign v_G1_2083_out0 = v_CARRY_2652_out0 || v_CARRY_2651_out0;
assign v_COUT_467_out0 = v_G1_2083_out0;
assign v__1373_out0 = { v__997_out0,v_S_731_out0 };
assign v_CIN_4972_out0 = v_COUT_467_out0;
assign v_RD_3161_out0 = v_CIN_4972_out0;
assign v_G1_4080_out0 = ((v_RD_3161_out0 && !v_RM_5852_out0) || (!v_RD_3161_out0) && v_RM_5852_out0);
assign v_G2_6325_out0 = v_RD_3161_out0 && v_RM_5852_out0;
assign v_CARRY_2662_out0 = v_G2_6325_out0;
assign v_S_4649_out0 = v_G1_4080_out0;
assign v_S_736_out0 = v_S_4649_out0;
assign v_G1_2088_out0 = v_CARRY_2662_out0 || v_CARRY_2661_out0;
assign v_COUT_472_out0 = v_G1_2088_out0;
assign v__900_out0 = { v__1373_out0,v_S_736_out0 };
assign v_CIN_4968_out0 = v_COUT_472_out0;
assign v_RD_3153_out0 = v_CIN_4968_out0;
assign v_G1_4072_out0 = ((v_RD_3153_out0 && !v_RM_5844_out0) || (!v_RD_3153_out0) && v_RM_5844_out0);
assign v_G2_6317_out0 = v_RD_3153_out0 && v_RM_5844_out0;
assign v_CARRY_2654_out0 = v_G2_6317_out0;
assign v_S_4641_out0 = v_G1_4072_out0;
assign v_S_732_out0 = v_S_4641_out0;
assign v_G1_2084_out0 = v_CARRY_2654_out0 || v_CARRY_2653_out0;
assign v_COUT_468_out0 = v_G1_2084_out0;
assign v__2229_out0 = { v__900_out0,v_S_732_out0 };
assign v_RM_1766_out0 = v_COUT_468_out0;
assign v_RM_5845_out0 = v_RM_1766_out0;
assign v_G1_4073_out0 = ((v_RD_3154_out0 && !v_RM_5845_out0) || (!v_RD_3154_out0) && v_RM_5845_out0);
assign v_G2_6318_out0 = v_RD_3154_out0 && v_RM_5845_out0;
assign v_CARRY_2655_out0 = v_G2_6318_out0;
assign v_S_4642_out0 = v_G1_4073_out0;
assign v_RM_5846_out0 = v_S_4642_out0;
assign v_G1_4074_out0 = ((v_RD_3155_out0 && !v_RM_5846_out0) || (!v_RD_3155_out0) && v_RM_5846_out0);
assign v_G2_6319_out0 = v_RD_3155_out0 && v_RM_5846_out0;
assign v_CARRY_2656_out0 = v_G2_6319_out0;
assign v_S_4643_out0 = v_G1_4074_out0;
assign v_S_733_out0 = v_S_4643_out0;
assign v_G1_2085_out0 = v_CARRY_2656_out0 || v_CARRY_2655_out0;
assign v_COUT_469_out0 = v_G1_2085_out0;
assign v__5252_out0 = { v__2229_out0,v_S_733_out0 };
assign v__5395_out0 = { v__5252_out0,v_COUT_469_out0 };
assign v_COUT_5380_out0 = v__5395_out0;
assign v_CIN_1161_out0 = v_COUT_5380_out0;
assign v__243_out0 = v_CIN_1161_out0[8:8];
assign v__881_out0 = v_CIN_1161_out0[6:6];
assign v__1064_out0 = v_CIN_1161_out0[3:3];
assign v__1083_out0 = v_CIN_1161_out0[15:15];
assign v__1234_out0 = v_CIN_1161_out0[0:0];
assign v__1502_out0 = v_CIN_1161_out0[9:9];
assign v__1518_out0 = v_CIN_1161_out0[2:2];
assign v__1544_out0 = v_CIN_1161_out0[7:7];
assign v__1877_out0 = v_CIN_1161_out0[1:1];
assign v__1895_out0 = v_CIN_1161_out0[10:10];
assign v__3354_out0 = v_CIN_1161_out0[11:11];
assign v__3770_out0 = v_CIN_1161_out0[12:12];
assign v__4296_out0 = v_CIN_1161_out0[13:13];
assign v__4329_out0 = v_CIN_1161_out0[14:14];
assign v__5290_out0 = v_CIN_1161_out0[5:5];
assign v__6638_out0 = v_CIN_1161_out0[4:4];
assign v_RM_1839_out0 = v__3770_out0;
assign v_RM_1840_out0 = v__4329_out0;
assign v_RM_1842_out0 = v__5290_out0;
assign v_RM_1843_out0 = v__6638_out0;
assign v_RM_1844_out0 = v__4296_out0;
assign v_RM_1845_out0 = v__1502_out0;
assign v_RM_1846_out0 = v__1895_out0;
assign v_RM_1847_out0 = v__1877_out0;
assign v_RM_1848_out0 = v__1064_out0;
assign v_RM_1849_out0 = v__881_out0;
assign v_RM_1850_out0 = v__1544_out0;
assign v_RM_1851_out0 = v__3354_out0;
assign v_RM_1852_out0 = v__243_out0;
assign v_RM_1853_out0 = v__1518_out0;
assign v_CIN_5044_out0 = v__1083_out0;
assign v_RM_6008_out0 = v__1234_out0;
assign v_RD_3310_out0 = v_CIN_5044_out0;
assign v_G1_4236_out0 = ((v_RD_3317_out0 && !v_RM_6008_out0) || (!v_RD_3317_out0) && v_RM_6008_out0);
assign v_RM_5996_out0 = v_RM_1839_out0;
assign v_RM_5998_out0 = v_RM_1840_out0;
assign v_RM_6002_out0 = v_RM_1842_out0;
assign v_RM_6004_out0 = v_RM_1843_out0;
assign v_RM_6006_out0 = v_RM_1844_out0;
assign v_RM_6009_out0 = v_RM_1845_out0;
assign v_RM_6011_out0 = v_RM_1846_out0;
assign v_RM_6013_out0 = v_RM_1847_out0;
assign v_RM_6015_out0 = v_RM_1848_out0;
assign v_RM_6017_out0 = v_RM_1849_out0;
assign v_RM_6019_out0 = v_RM_1850_out0;
assign v_RM_6021_out0 = v_RM_1851_out0;
assign v_RM_6023_out0 = v_RM_1852_out0;
assign v_RM_6025_out0 = v_RM_1853_out0;
assign v_G2_6481_out0 = v_RD_3317_out0 && v_RM_6008_out0;
assign v_CARRY_2818_out0 = v_G2_6481_out0;
assign v_G1_4224_out0 = ((v_RD_3305_out0 && !v_RM_5996_out0) || (!v_RD_3305_out0) && v_RM_5996_out0);
assign v_G1_4226_out0 = ((v_RD_3307_out0 && !v_RM_5998_out0) || (!v_RD_3307_out0) && v_RM_5998_out0);
assign v_G1_4230_out0 = ((v_RD_3311_out0 && !v_RM_6002_out0) || (!v_RD_3311_out0) && v_RM_6002_out0);
assign v_G1_4232_out0 = ((v_RD_3313_out0 && !v_RM_6004_out0) || (!v_RD_3313_out0) && v_RM_6004_out0);
assign v_G1_4234_out0 = ((v_RD_3315_out0 && !v_RM_6006_out0) || (!v_RD_3315_out0) && v_RM_6006_out0);
assign v_G1_4237_out0 = ((v_RD_3318_out0 && !v_RM_6009_out0) || (!v_RD_3318_out0) && v_RM_6009_out0);
assign v_G1_4239_out0 = ((v_RD_3320_out0 && !v_RM_6011_out0) || (!v_RD_3320_out0) && v_RM_6011_out0);
assign v_G1_4241_out0 = ((v_RD_3322_out0 && !v_RM_6013_out0) || (!v_RD_3322_out0) && v_RM_6013_out0);
assign v_G1_4243_out0 = ((v_RD_3324_out0 && !v_RM_6015_out0) || (!v_RD_3324_out0) && v_RM_6015_out0);
assign v_G1_4245_out0 = ((v_RD_3326_out0 && !v_RM_6017_out0) || (!v_RD_3326_out0) && v_RM_6017_out0);
assign v_G1_4247_out0 = ((v_RD_3328_out0 && !v_RM_6019_out0) || (!v_RD_3328_out0) && v_RM_6019_out0);
assign v_G1_4249_out0 = ((v_RD_3330_out0 && !v_RM_6021_out0) || (!v_RD_3330_out0) && v_RM_6021_out0);
assign v_G1_4251_out0 = ((v_RD_3332_out0 && !v_RM_6023_out0) || (!v_RD_3332_out0) && v_RM_6023_out0);
assign v_G1_4253_out0 = ((v_RD_3334_out0 && !v_RM_6025_out0) || (!v_RD_3334_out0) && v_RM_6025_out0);
assign v_S_4805_out0 = v_G1_4236_out0;
assign v_G2_6469_out0 = v_RD_3305_out0 && v_RM_5996_out0;
assign v_G2_6471_out0 = v_RD_3307_out0 && v_RM_5998_out0;
assign v_G2_6475_out0 = v_RD_3311_out0 && v_RM_6002_out0;
assign v_G2_6477_out0 = v_RD_3313_out0 && v_RM_6004_out0;
assign v_G2_6479_out0 = v_RD_3315_out0 && v_RM_6006_out0;
assign v_G2_6482_out0 = v_RD_3318_out0 && v_RM_6009_out0;
assign v_G2_6484_out0 = v_RD_3320_out0 && v_RM_6011_out0;
assign v_G2_6486_out0 = v_RD_3322_out0 && v_RM_6013_out0;
assign v_G2_6488_out0 = v_RD_3324_out0 && v_RM_6015_out0;
assign v_G2_6490_out0 = v_RD_3326_out0 && v_RM_6017_out0;
assign v_G2_6492_out0 = v_RD_3328_out0 && v_RM_6019_out0;
assign v_G2_6494_out0 = v_RD_3330_out0 && v_RM_6021_out0;
assign v_G2_6496_out0 = v_RD_3332_out0 && v_RM_6023_out0;
assign v_G2_6498_out0 = v_RD_3334_out0 && v_RM_6025_out0;
assign v_S_2292_out0 = v_S_4805_out0;
assign v_CARRY_2806_out0 = v_G2_6469_out0;
assign v_CARRY_2808_out0 = v_G2_6471_out0;
assign v_CARRY_2812_out0 = v_G2_6475_out0;
assign v_CARRY_2814_out0 = v_G2_6477_out0;
assign v_CARRY_2816_out0 = v_G2_6479_out0;
assign v_CARRY_2819_out0 = v_G2_6482_out0;
assign v_CARRY_2821_out0 = v_G2_6484_out0;
assign v_CARRY_2823_out0 = v_G2_6486_out0;
assign v_CARRY_2825_out0 = v_G2_6488_out0;
assign v_CARRY_2827_out0 = v_G2_6490_out0;
assign v_CARRY_2829_out0 = v_G2_6492_out0;
assign v_CARRY_2831_out0 = v_G2_6494_out0;
assign v_CARRY_2833_out0 = v_G2_6496_out0;
assign v_CARRY_2835_out0 = v_G2_6498_out0;
assign v_S_4793_out0 = v_G1_4224_out0;
assign v_S_4795_out0 = v_G1_4226_out0;
assign v_S_4799_out0 = v_G1_4230_out0;
assign v_S_4801_out0 = v_G1_4232_out0;
assign v_S_4803_out0 = v_G1_4234_out0;
assign v_S_4806_out0 = v_G1_4237_out0;
assign v_S_4808_out0 = v_G1_4239_out0;
assign v_S_4810_out0 = v_G1_4241_out0;
assign v_S_4812_out0 = v_G1_4243_out0;
assign v_S_4814_out0 = v_G1_4245_out0;
assign v_S_4816_out0 = v_G1_4247_out0;
assign v_S_4818_out0 = v_G1_4249_out0;
assign v_S_4820_out0 = v_G1_4251_out0;
assign v_S_4822_out0 = v_G1_4253_out0;
assign v_CIN_5050_out0 = v_CARRY_2818_out0;
assign v_RD_3323_out0 = v_CIN_5050_out0;
assign v__5303_out0 = { v__24_out0,v_S_2292_out0 };
assign v_RM_5997_out0 = v_S_4793_out0;
assign v_RM_5999_out0 = v_S_4795_out0;
assign v_RM_6003_out0 = v_S_4799_out0;
assign v_RM_6005_out0 = v_S_4801_out0;
assign v_RM_6007_out0 = v_S_4803_out0;
assign v_RM_6010_out0 = v_S_4806_out0;
assign v_RM_6012_out0 = v_S_4808_out0;
assign v_RM_6014_out0 = v_S_4810_out0;
assign v_RM_6016_out0 = v_S_4812_out0;
assign v_RM_6018_out0 = v_S_4814_out0;
assign v_RM_6020_out0 = v_S_4816_out0;
assign v_RM_6022_out0 = v_S_4818_out0;
assign v_RM_6024_out0 = v_S_4820_out0;
assign v_RM_6026_out0 = v_S_4822_out0;
assign v_G1_4242_out0 = ((v_RD_3323_out0 && !v_RM_6014_out0) || (!v_RD_3323_out0) && v_RM_6014_out0);
assign v_G2_6487_out0 = v_RD_3323_out0 && v_RM_6014_out0;
assign v_CARRY_2824_out0 = v_G2_6487_out0;
assign v_S_4811_out0 = v_G1_4242_out0;
assign v_S_814_out0 = v_S_4811_out0;
assign v_G1_2166_out0 = v_CARRY_2824_out0 || v_CARRY_2823_out0;
assign v_COUT_550_out0 = v_G1_2166_out0;
assign v_CIN_5056_out0 = v_COUT_550_out0;
assign v_RD_3335_out0 = v_CIN_5056_out0;
assign v_G1_4254_out0 = ((v_RD_3335_out0 && !v_RM_6026_out0) || (!v_RD_3335_out0) && v_RM_6026_out0);
assign v_G2_6499_out0 = v_RD_3335_out0 && v_RM_6026_out0;
assign v_CARRY_2836_out0 = v_G2_6499_out0;
assign v_S_4823_out0 = v_G1_4254_out0;
assign v_S_820_out0 = v_S_4823_out0;
assign v_G1_2172_out0 = v_CARRY_2836_out0 || v_CARRY_2835_out0;
assign v_COUT_556_out0 = v_G1_2172_out0;
assign v__2349_out0 = { v_S_814_out0,v_S_820_out0 };
assign v_CIN_5051_out0 = v_COUT_556_out0;
assign v_RD_3325_out0 = v_CIN_5051_out0;
assign v_G1_4244_out0 = ((v_RD_3325_out0 && !v_RM_6016_out0) || (!v_RD_3325_out0) && v_RM_6016_out0);
assign v_G2_6489_out0 = v_RD_3325_out0 && v_RM_6016_out0;
assign v_CARRY_2826_out0 = v_G2_6489_out0;
assign v_S_4813_out0 = v_G1_4244_out0;
assign v_S_815_out0 = v_S_4813_out0;
assign v_G1_2167_out0 = v_CARRY_2826_out0 || v_CARRY_2825_out0;
assign v_COUT_551_out0 = v_G1_2167_out0;
assign v__1258_out0 = { v__2349_out0,v_S_815_out0 };
assign v_CIN_5046_out0 = v_COUT_551_out0;
assign v_RD_3314_out0 = v_CIN_5046_out0;
assign v_G1_4233_out0 = ((v_RD_3314_out0 && !v_RM_6005_out0) || (!v_RD_3314_out0) && v_RM_6005_out0);
assign v_G2_6478_out0 = v_RD_3314_out0 && v_RM_6005_out0;
assign v_CARRY_2815_out0 = v_G2_6478_out0;
assign v_S_4802_out0 = v_G1_4233_out0;
assign v_S_810_out0 = v_S_4802_out0;
assign v_G1_2162_out0 = v_CARRY_2815_out0 || v_CARRY_2814_out0;
assign v_COUT_546_out0 = v_G1_2162_out0;
assign v__3466_out0 = { v__1258_out0,v_S_810_out0 };
assign v_CIN_5045_out0 = v_COUT_546_out0;
assign v_RD_3312_out0 = v_CIN_5045_out0;
assign v_G1_4231_out0 = ((v_RD_3312_out0 && !v_RM_6003_out0) || (!v_RD_3312_out0) && v_RM_6003_out0);
assign v_G2_6476_out0 = v_RD_3312_out0 && v_RM_6003_out0;
assign v_CARRY_2813_out0 = v_G2_6476_out0;
assign v_S_4800_out0 = v_G1_4231_out0;
assign v_S_809_out0 = v_S_4800_out0;
assign v_G1_2161_out0 = v_CARRY_2813_out0 || v_CARRY_2812_out0;
assign v_COUT_545_out0 = v_G1_2161_out0;
assign v__6676_out0 = { v__3466_out0,v_S_809_out0 };
assign v_CIN_5052_out0 = v_COUT_545_out0;
assign v_RD_3327_out0 = v_CIN_5052_out0;
assign v_G1_4246_out0 = ((v_RD_3327_out0 && !v_RM_6018_out0) || (!v_RD_3327_out0) && v_RM_6018_out0);
assign v_G2_6491_out0 = v_RD_3327_out0 && v_RM_6018_out0;
assign v_CARRY_2828_out0 = v_G2_6491_out0;
assign v_S_4815_out0 = v_G1_4246_out0;
assign v_S_816_out0 = v_S_4815_out0;
assign v_G1_2168_out0 = v_CARRY_2828_out0 || v_CARRY_2827_out0;
assign v_COUT_552_out0 = v_G1_2168_out0;
assign v__1624_out0 = { v__6676_out0,v_S_816_out0 };
assign v_CIN_5053_out0 = v_COUT_552_out0;
assign v_RD_3329_out0 = v_CIN_5053_out0;
assign v_G1_4248_out0 = ((v_RD_3329_out0 && !v_RM_6020_out0) || (!v_RD_3329_out0) && v_RM_6020_out0);
assign v_G2_6493_out0 = v_RD_3329_out0 && v_RM_6020_out0;
assign v_CARRY_2830_out0 = v_G2_6493_out0;
assign v_S_4817_out0 = v_G1_4248_out0;
assign v_S_817_out0 = v_S_4817_out0;
assign v_G1_2169_out0 = v_CARRY_2830_out0 || v_CARRY_2829_out0;
assign v_COUT_553_out0 = v_G1_2169_out0;
assign v__3521_out0 = { v__1624_out0,v_S_817_out0 };
assign v_CIN_5055_out0 = v_COUT_553_out0;
assign v_RD_3333_out0 = v_CIN_5055_out0;
assign v_G1_4252_out0 = ((v_RD_3333_out0 && !v_RM_6024_out0) || (!v_RD_3333_out0) && v_RM_6024_out0);
assign v_G2_6497_out0 = v_RD_3333_out0 && v_RM_6024_out0;
assign v_CARRY_2834_out0 = v_G2_6497_out0;
assign v_S_4821_out0 = v_G1_4252_out0;
assign v_S_819_out0 = v_S_4821_out0;
assign v_G1_2171_out0 = v_CARRY_2834_out0 || v_CARRY_2833_out0;
assign v_COUT_555_out0 = v_G1_2171_out0;
assign v__2332_out0 = { v__3521_out0,v_S_819_out0 };
assign v_CIN_5048_out0 = v_COUT_555_out0;
assign v_RD_3319_out0 = v_CIN_5048_out0;
assign v_G1_4238_out0 = ((v_RD_3319_out0 && !v_RM_6010_out0) || (!v_RD_3319_out0) && v_RM_6010_out0);
assign v_G2_6483_out0 = v_RD_3319_out0 && v_RM_6010_out0;
assign v_CARRY_2820_out0 = v_G2_6483_out0;
assign v_S_4807_out0 = v_G1_4238_out0;
assign v_S_812_out0 = v_S_4807_out0;
assign v_G1_2164_out0 = v_CARRY_2820_out0 || v_CARRY_2819_out0;
assign v_COUT_548_out0 = v_G1_2164_out0;
assign v__3414_out0 = { v__2332_out0,v_S_812_out0 };
assign v_CIN_5049_out0 = v_COUT_548_out0;
assign v_RD_3321_out0 = v_CIN_5049_out0;
assign v_G1_4240_out0 = ((v_RD_3321_out0 && !v_RM_6012_out0) || (!v_RD_3321_out0) && v_RM_6012_out0);
assign v_G2_6485_out0 = v_RD_3321_out0 && v_RM_6012_out0;
assign v_CARRY_2822_out0 = v_G2_6485_out0;
assign v_S_4809_out0 = v_G1_4240_out0;
assign v_S_813_out0 = v_S_4809_out0;
assign v_G1_2165_out0 = v_CARRY_2822_out0 || v_CARRY_2821_out0;
assign v_COUT_549_out0 = v_G1_2165_out0;
assign v__2858_out0 = { v__3414_out0,v_S_813_out0 };
assign v_CIN_5054_out0 = v_COUT_549_out0;
assign v_RD_3331_out0 = v_CIN_5054_out0;
assign v_G1_4250_out0 = ((v_RD_3331_out0 && !v_RM_6022_out0) || (!v_RD_3331_out0) && v_RM_6022_out0);
assign v_G2_6495_out0 = v_RD_3331_out0 && v_RM_6022_out0;
assign v_CARRY_2832_out0 = v_G2_6495_out0;
assign v_S_4819_out0 = v_G1_4250_out0;
assign v_S_818_out0 = v_S_4819_out0;
assign v_G1_2170_out0 = v_CARRY_2832_out0 || v_CARRY_2831_out0;
assign v_COUT_554_out0 = v_G1_2170_out0;
assign v__1002_out0 = { v__2858_out0,v_S_818_out0 };
assign v_CIN_5042_out0 = v_COUT_554_out0;
assign v_RD_3306_out0 = v_CIN_5042_out0;
assign v_G1_4225_out0 = ((v_RD_3306_out0 && !v_RM_5997_out0) || (!v_RD_3306_out0) && v_RM_5997_out0);
assign v_G2_6470_out0 = v_RD_3306_out0 && v_RM_5997_out0;
assign v_CARRY_2807_out0 = v_G2_6470_out0;
assign v_S_4794_out0 = v_G1_4225_out0;
assign v_S_806_out0 = v_S_4794_out0;
assign v_G1_2158_out0 = v_CARRY_2807_out0 || v_CARRY_2806_out0;
assign v_COUT_542_out0 = v_G1_2158_out0;
assign v__1378_out0 = { v__1002_out0,v_S_806_out0 };
assign v_CIN_5047_out0 = v_COUT_542_out0;
assign v_RD_3316_out0 = v_CIN_5047_out0;
assign v_G1_4235_out0 = ((v_RD_3316_out0 && !v_RM_6007_out0) || (!v_RD_3316_out0) && v_RM_6007_out0);
assign v_G2_6480_out0 = v_RD_3316_out0 && v_RM_6007_out0;
assign v_CARRY_2817_out0 = v_G2_6480_out0;
assign v_S_4804_out0 = v_G1_4235_out0;
assign v_S_811_out0 = v_S_4804_out0;
assign v_G1_2163_out0 = v_CARRY_2817_out0 || v_CARRY_2816_out0;
assign v_COUT_547_out0 = v_G1_2163_out0;
assign v__905_out0 = { v__1378_out0,v_S_811_out0 };
assign v_CIN_5043_out0 = v_COUT_547_out0;
assign v_RD_3308_out0 = v_CIN_5043_out0;
assign v_G1_4227_out0 = ((v_RD_3308_out0 && !v_RM_5999_out0) || (!v_RD_3308_out0) && v_RM_5999_out0);
assign v_G2_6472_out0 = v_RD_3308_out0 && v_RM_5999_out0;
assign v_CARRY_2809_out0 = v_G2_6472_out0;
assign v_S_4796_out0 = v_G1_4227_out0;
assign v_S_807_out0 = v_S_4796_out0;
assign v_G1_2159_out0 = v_CARRY_2809_out0 || v_CARRY_2808_out0;
assign v_COUT_543_out0 = v_G1_2159_out0;
assign v__2234_out0 = { v__905_out0,v_S_807_out0 };
assign v_RM_1841_out0 = v_COUT_543_out0;
assign v_RM_6000_out0 = v_RM_1841_out0;
assign v_G1_4228_out0 = ((v_RD_3309_out0 && !v_RM_6000_out0) || (!v_RD_3309_out0) && v_RM_6000_out0);
assign v_G2_6473_out0 = v_RD_3309_out0 && v_RM_6000_out0;
assign v_CARRY_2810_out0 = v_G2_6473_out0;
assign v_S_4797_out0 = v_G1_4228_out0;
assign v_RM_6001_out0 = v_S_4797_out0;
assign v_G1_4229_out0 = ((v_RD_3310_out0 && !v_RM_6001_out0) || (!v_RD_3310_out0) && v_RM_6001_out0);
assign v_G2_6474_out0 = v_RD_3310_out0 && v_RM_6001_out0;
assign v_CARRY_2811_out0 = v_G2_6474_out0;
assign v_S_4798_out0 = v_G1_4229_out0;
assign v_S_808_out0 = v_S_4798_out0;
assign v_G1_2160_out0 = v_CARRY_2811_out0 || v_CARRY_2810_out0;
assign v_COUT_544_out0 = v_G1_2160_out0;
assign v__5257_out0 = { v__2234_out0,v_S_808_out0 };
assign v__5400_out0 = { v__5257_out0,v_COUT_544_out0 };
assign v_COUT_5385_out0 = v__5400_out0;
assign v_CIN_1152_out0 = v_COUT_5385_out0;
assign v__234_out0 = v_CIN_1152_out0[8:8];
assign v__872_out0 = v_CIN_1152_out0[6:6];
assign v__1055_out0 = v_CIN_1152_out0[3:3];
assign v__1074_out0 = v_CIN_1152_out0[15:15];
assign v__1225_out0 = v_CIN_1152_out0[0:0];
assign v__1493_out0 = v_CIN_1152_out0[9:9];
assign v__1509_out0 = v_CIN_1152_out0[2:2];
assign v__1535_out0 = v_CIN_1152_out0[7:7];
assign v__1868_out0 = v_CIN_1152_out0[1:1];
assign v__1886_out0 = v_CIN_1152_out0[10:10];
assign v__3345_out0 = v_CIN_1152_out0[11:11];
assign v__3761_out0 = v_CIN_1152_out0[12:12];
assign v__4287_out0 = v_CIN_1152_out0[13:13];
assign v__4320_out0 = v_CIN_1152_out0[14:14];
assign v__5281_out0 = v_CIN_1152_out0[5:5];
assign v__6629_out0 = v_CIN_1152_out0[4:4];
assign v_RM_1704_out0 = v__3761_out0;
assign v_RM_1705_out0 = v__4320_out0;
assign v_RM_1707_out0 = v__5281_out0;
assign v_RM_1708_out0 = v__6629_out0;
assign v_RM_1709_out0 = v__4287_out0;
assign v_RM_1710_out0 = v__1493_out0;
assign v_RM_1711_out0 = v__1886_out0;
assign v_RM_1712_out0 = v__1868_out0;
assign v_RM_1713_out0 = v__1055_out0;
assign v_RM_1714_out0 = v__872_out0;
assign v_RM_1715_out0 = v__1535_out0;
assign v_RM_1716_out0 = v__3345_out0;
assign v_RM_1717_out0 = v__234_out0;
assign v_RM_1718_out0 = v__1509_out0;
assign v_CIN_4909_out0 = v__1074_out0;
assign v_RM_5729_out0 = v__1225_out0;
assign v_RD_3031_out0 = v_CIN_4909_out0;
assign v_G1_3957_out0 = ((v_RD_3038_out0 && !v_RM_5729_out0) || (!v_RD_3038_out0) && v_RM_5729_out0);
assign v_RM_5717_out0 = v_RM_1704_out0;
assign v_RM_5719_out0 = v_RM_1705_out0;
assign v_RM_5723_out0 = v_RM_1707_out0;
assign v_RM_5725_out0 = v_RM_1708_out0;
assign v_RM_5727_out0 = v_RM_1709_out0;
assign v_RM_5730_out0 = v_RM_1710_out0;
assign v_RM_5732_out0 = v_RM_1711_out0;
assign v_RM_5734_out0 = v_RM_1712_out0;
assign v_RM_5736_out0 = v_RM_1713_out0;
assign v_RM_5738_out0 = v_RM_1714_out0;
assign v_RM_5740_out0 = v_RM_1715_out0;
assign v_RM_5742_out0 = v_RM_1716_out0;
assign v_RM_5744_out0 = v_RM_1717_out0;
assign v_RM_5746_out0 = v_RM_1718_out0;
assign v_G2_6202_out0 = v_RD_3038_out0 && v_RM_5729_out0;
assign v_CARRY_2539_out0 = v_G2_6202_out0;
assign v_G1_3945_out0 = ((v_RD_3026_out0 && !v_RM_5717_out0) || (!v_RD_3026_out0) && v_RM_5717_out0);
assign v_G1_3947_out0 = ((v_RD_3028_out0 && !v_RM_5719_out0) || (!v_RD_3028_out0) && v_RM_5719_out0);
assign v_G1_3951_out0 = ((v_RD_3032_out0 && !v_RM_5723_out0) || (!v_RD_3032_out0) && v_RM_5723_out0);
assign v_G1_3953_out0 = ((v_RD_3034_out0 && !v_RM_5725_out0) || (!v_RD_3034_out0) && v_RM_5725_out0);
assign v_G1_3955_out0 = ((v_RD_3036_out0 && !v_RM_5727_out0) || (!v_RD_3036_out0) && v_RM_5727_out0);
assign v_G1_3958_out0 = ((v_RD_3039_out0 && !v_RM_5730_out0) || (!v_RD_3039_out0) && v_RM_5730_out0);
assign v_G1_3960_out0 = ((v_RD_3041_out0 && !v_RM_5732_out0) || (!v_RD_3041_out0) && v_RM_5732_out0);
assign v_G1_3962_out0 = ((v_RD_3043_out0 && !v_RM_5734_out0) || (!v_RD_3043_out0) && v_RM_5734_out0);
assign v_G1_3964_out0 = ((v_RD_3045_out0 && !v_RM_5736_out0) || (!v_RD_3045_out0) && v_RM_5736_out0);
assign v_G1_3966_out0 = ((v_RD_3047_out0 && !v_RM_5738_out0) || (!v_RD_3047_out0) && v_RM_5738_out0);
assign v_G1_3968_out0 = ((v_RD_3049_out0 && !v_RM_5740_out0) || (!v_RD_3049_out0) && v_RM_5740_out0);
assign v_G1_3970_out0 = ((v_RD_3051_out0 && !v_RM_5742_out0) || (!v_RD_3051_out0) && v_RM_5742_out0);
assign v_G1_3972_out0 = ((v_RD_3053_out0 && !v_RM_5744_out0) || (!v_RD_3053_out0) && v_RM_5744_out0);
assign v_G1_3974_out0 = ((v_RD_3055_out0 && !v_RM_5746_out0) || (!v_RD_3055_out0) && v_RM_5746_out0);
assign v_S_4526_out0 = v_G1_3957_out0;
assign v_G2_6190_out0 = v_RD_3026_out0 && v_RM_5717_out0;
assign v_G2_6192_out0 = v_RD_3028_out0 && v_RM_5719_out0;
assign v_G2_6196_out0 = v_RD_3032_out0 && v_RM_5723_out0;
assign v_G2_6198_out0 = v_RD_3034_out0 && v_RM_5725_out0;
assign v_G2_6200_out0 = v_RD_3036_out0 && v_RM_5727_out0;
assign v_G2_6203_out0 = v_RD_3039_out0 && v_RM_5730_out0;
assign v_G2_6205_out0 = v_RD_3041_out0 && v_RM_5732_out0;
assign v_G2_6207_out0 = v_RD_3043_out0 && v_RM_5734_out0;
assign v_G2_6209_out0 = v_RD_3045_out0 && v_RM_5736_out0;
assign v_G2_6211_out0 = v_RD_3047_out0 && v_RM_5738_out0;
assign v_G2_6213_out0 = v_RD_3049_out0 && v_RM_5740_out0;
assign v_G2_6215_out0 = v_RD_3051_out0 && v_RM_5742_out0;
assign v_G2_6217_out0 = v_RD_3053_out0 && v_RM_5744_out0;
assign v_G2_6219_out0 = v_RD_3055_out0 && v_RM_5746_out0;
assign v_S_2283_out0 = v_S_4526_out0;
assign v_CARRY_2527_out0 = v_G2_6190_out0;
assign v_CARRY_2529_out0 = v_G2_6192_out0;
assign v_CARRY_2533_out0 = v_G2_6196_out0;
assign v_CARRY_2535_out0 = v_G2_6198_out0;
assign v_CARRY_2537_out0 = v_G2_6200_out0;
assign v_CARRY_2540_out0 = v_G2_6203_out0;
assign v_CARRY_2542_out0 = v_G2_6205_out0;
assign v_CARRY_2544_out0 = v_G2_6207_out0;
assign v_CARRY_2546_out0 = v_G2_6209_out0;
assign v_CARRY_2548_out0 = v_G2_6211_out0;
assign v_CARRY_2550_out0 = v_G2_6213_out0;
assign v_CARRY_2552_out0 = v_G2_6215_out0;
assign v_CARRY_2554_out0 = v_G2_6217_out0;
assign v_CARRY_2556_out0 = v_G2_6219_out0;
assign v_S_4514_out0 = v_G1_3945_out0;
assign v_S_4516_out0 = v_G1_3947_out0;
assign v_S_4520_out0 = v_G1_3951_out0;
assign v_S_4522_out0 = v_G1_3953_out0;
assign v_S_4524_out0 = v_G1_3955_out0;
assign v_S_4527_out0 = v_G1_3958_out0;
assign v_S_4529_out0 = v_G1_3960_out0;
assign v_S_4531_out0 = v_G1_3962_out0;
assign v_S_4533_out0 = v_G1_3964_out0;
assign v_S_4535_out0 = v_G1_3966_out0;
assign v_S_4537_out0 = v_G1_3968_out0;
assign v_S_4539_out0 = v_G1_3970_out0;
assign v_S_4541_out0 = v_G1_3972_out0;
assign v_S_4543_out0 = v_G1_3974_out0;
assign v_CIN_4915_out0 = v_CARRY_2539_out0;
assign v__1068_out0 = { v__5303_out0,v_S_2283_out0 };
assign v_RD_3044_out0 = v_CIN_4915_out0;
assign v_RM_5718_out0 = v_S_4514_out0;
assign v_RM_5720_out0 = v_S_4516_out0;
assign v_RM_5724_out0 = v_S_4520_out0;
assign v_RM_5726_out0 = v_S_4522_out0;
assign v_RM_5728_out0 = v_S_4524_out0;
assign v_RM_5731_out0 = v_S_4527_out0;
assign v_RM_5733_out0 = v_S_4529_out0;
assign v_RM_5735_out0 = v_S_4531_out0;
assign v_RM_5737_out0 = v_S_4533_out0;
assign v_RM_5739_out0 = v_S_4535_out0;
assign v_RM_5741_out0 = v_S_4537_out0;
assign v_RM_5743_out0 = v_S_4539_out0;
assign v_RM_5745_out0 = v_S_4541_out0;
assign v_RM_5747_out0 = v_S_4543_out0;
assign v_G1_3963_out0 = ((v_RD_3044_out0 && !v_RM_5735_out0) || (!v_RD_3044_out0) && v_RM_5735_out0);
assign v_G2_6208_out0 = v_RD_3044_out0 && v_RM_5735_out0;
assign v_CARRY_2545_out0 = v_G2_6208_out0;
assign v_S_4532_out0 = v_G1_3963_out0;
assign v_S_679_out0 = v_S_4532_out0;
assign v_G1_2031_out0 = v_CARRY_2545_out0 || v_CARRY_2544_out0;
assign v_COUT_415_out0 = v_G1_2031_out0;
assign v_CIN_4921_out0 = v_COUT_415_out0;
assign v_RD_3056_out0 = v_CIN_4921_out0;
assign v_G1_3975_out0 = ((v_RD_3056_out0 && !v_RM_5747_out0) || (!v_RD_3056_out0) && v_RM_5747_out0);
assign v_G2_6220_out0 = v_RD_3056_out0 && v_RM_5747_out0;
assign v_CARRY_2557_out0 = v_G2_6220_out0;
assign v_S_4544_out0 = v_G1_3975_out0;
assign v_S_685_out0 = v_S_4544_out0;
assign v_G1_2037_out0 = v_CARRY_2557_out0 || v_CARRY_2556_out0;
assign v_COUT_421_out0 = v_G1_2037_out0;
assign v__2340_out0 = { v_S_679_out0,v_S_685_out0 };
assign v_CIN_4916_out0 = v_COUT_421_out0;
assign v_RD_3046_out0 = v_CIN_4916_out0;
assign v_G1_3965_out0 = ((v_RD_3046_out0 && !v_RM_5737_out0) || (!v_RD_3046_out0) && v_RM_5737_out0);
assign v_G2_6210_out0 = v_RD_3046_out0 && v_RM_5737_out0;
assign v_CARRY_2547_out0 = v_G2_6210_out0;
assign v_S_4534_out0 = v_G1_3965_out0;
assign v_S_680_out0 = v_S_4534_out0;
assign v_G1_2032_out0 = v_CARRY_2547_out0 || v_CARRY_2546_out0;
assign v_COUT_416_out0 = v_G1_2032_out0;
assign v__1249_out0 = { v__2340_out0,v_S_680_out0 };
assign v_CIN_4911_out0 = v_COUT_416_out0;
assign v_RD_3035_out0 = v_CIN_4911_out0;
assign v_G1_3954_out0 = ((v_RD_3035_out0 && !v_RM_5726_out0) || (!v_RD_3035_out0) && v_RM_5726_out0);
assign v_G2_6199_out0 = v_RD_3035_out0 && v_RM_5726_out0;
assign v_CARRY_2536_out0 = v_G2_6199_out0;
assign v_S_4523_out0 = v_G1_3954_out0;
assign v_S_675_out0 = v_S_4523_out0;
assign v_G1_2027_out0 = v_CARRY_2536_out0 || v_CARRY_2535_out0;
assign v_COUT_411_out0 = v_G1_2027_out0;
assign v__3457_out0 = { v__1249_out0,v_S_675_out0 };
assign v_CIN_4910_out0 = v_COUT_411_out0;
assign v_RD_3033_out0 = v_CIN_4910_out0;
assign v_G1_3952_out0 = ((v_RD_3033_out0 && !v_RM_5724_out0) || (!v_RD_3033_out0) && v_RM_5724_out0);
assign v_G2_6197_out0 = v_RD_3033_out0 && v_RM_5724_out0;
assign v_CARRY_2534_out0 = v_G2_6197_out0;
assign v_S_4521_out0 = v_G1_3952_out0;
assign v_S_674_out0 = v_S_4521_out0;
assign v_G1_2026_out0 = v_CARRY_2534_out0 || v_CARRY_2533_out0;
assign v_COUT_410_out0 = v_G1_2026_out0;
assign v__6667_out0 = { v__3457_out0,v_S_674_out0 };
assign v_CIN_4917_out0 = v_COUT_410_out0;
assign v_RD_3048_out0 = v_CIN_4917_out0;
assign v_G1_3967_out0 = ((v_RD_3048_out0 && !v_RM_5739_out0) || (!v_RD_3048_out0) && v_RM_5739_out0);
assign v_G2_6212_out0 = v_RD_3048_out0 && v_RM_5739_out0;
assign v_CARRY_2549_out0 = v_G2_6212_out0;
assign v_S_4536_out0 = v_G1_3967_out0;
assign v_S_681_out0 = v_S_4536_out0;
assign v_G1_2033_out0 = v_CARRY_2549_out0 || v_CARRY_2548_out0;
assign v_COUT_417_out0 = v_G1_2033_out0;
assign v__1615_out0 = { v__6667_out0,v_S_681_out0 };
assign v_CIN_4918_out0 = v_COUT_417_out0;
assign v_RD_3050_out0 = v_CIN_4918_out0;
assign v_G1_3969_out0 = ((v_RD_3050_out0 && !v_RM_5741_out0) || (!v_RD_3050_out0) && v_RM_5741_out0);
assign v_G2_6214_out0 = v_RD_3050_out0 && v_RM_5741_out0;
assign v_CARRY_2551_out0 = v_G2_6214_out0;
assign v_S_4538_out0 = v_G1_3969_out0;
assign v_S_682_out0 = v_S_4538_out0;
assign v_G1_2034_out0 = v_CARRY_2551_out0 || v_CARRY_2550_out0;
assign v_COUT_418_out0 = v_G1_2034_out0;
assign v__3512_out0 = { v__1615_out0,v_S_682_out0 };
assign v_CIN_4920_out0 = v_COUT_418_out0;
assign v_RD_3054_out0 = v_CIN_4920_out0;
assign v_G1_3973_out0 = ((v_RD_3054_out0 && !v_RM_5745_out0) || (!v_RD_3054_out0) && v_RM_5745_out0);
assign v_G2_6218_out0 = v_RD_3054_out0 && v_RM_5745_out0;
assign v_CARRY_2555_out0 = v_G2_6218_out0;
assign v_S_4542_out0 = v_G1_3973_out0;
assign v_S_684_out0 = v_S_4542_out0;
assign v_G1_2036_out0 = v_CARRY_2555_out0 || v_CARRY_2554_out0;
assign v_COUT_420_out0 = v_G1_2036_out0;
assign v__2323_out0 = { v__3512_out0,v_S_684_out0 };
assign v_CIN_4913_out0 = v_COUT_420_out0;
assign v_RD_3040_out0 = v_CIN_4913_out0;
assign v_G1_3959_out0 = ((v_RD_3040_out0 && !v_RM_5731_out0) || (!v_RD_3040_out0) && v_RM_5731_out0);
assign v_G2_6204_out0 = v_RD_3040_out0 && v_RM_5731_out0;
assign v_CARRY_2541_out0 = v_G2_6204_out0;
assign v_S_4528_out0 = v_G1_3959_out0;
assign v_S_677_out0 = v_S_4528_out0;
assign v_G1_2029_out0 = v_CARRY_2541_out0 || v_CARRY_2540_out0;
assign v_COUT_413_out0 = v_G1_2029_out0;
assign v__3405_out0 = { v__2323_out0,v_S_677_out0 };
assign v_CIN_4914_out0 = v_COUT_413_out0;
assign v_RD_3042_out0 = v_CIN_4914_out0;
assign v_G1_3961_out0 = ((v_RD_3042_out0 && !v_RM_5733_out0) || (!v_RD_3042_out0) && v_RM_5733_out0);
assign v_G2_6206_out0 = v_RD_3042_out0 && v_RM_5733_out0;
assign v_CARRY_2543_out0 = v_G2_6206_out0;
assign v_S_4530_out0 = v_G1_3961_out0;
assign v_S_678_out0 = v_S_4530_out0;
assign v_G1_2030_out0 = v_CARRY_2543_out0 || v_CARRY_2542_out0;
assign v_COUT_414_out0 = v_G1_2030_out0;
assign v__2849_out0 = { v__3405_out0,v_S_678_out0 };
assign v_CIN_4919_out0 = v_COUT_414_out0;
assign v_RD_3052_out0 = v_CIN_4919_out0;
assign v_G1_3971_out0 = ((v_RD_3052_out0 && !v_RM_5743_out0) || (!v_RD_3052_out0) && v_RM_5743_out0);
assign v_G2_6216_out0 = v_RD_3052_out0 && v_RM_5743_out0;
assign v_CARRY_2553_out0 = v_G2_6216_out0;
assign v_S_4540_out0 = v_G1_3971_out0;
assign v_S_683_out0 = v_S_4540_out0;
assign v_G1_2035_out0 = v_CARRY_2553_out0 || v_CARRY_2552_out0;
assign v_COUT_419_out0 = v_G1_2035_out0;
assign v__993_out0 = { v__2849_out0,v_S_683_out0 };
assign v_CIN_4907_out0 = v_COUT_419_out0;
assign v_RD_3027_out0 = v_CIN_4907_out0;
assign v_G1_3946_out0 = ((v_RD_3027_out0 && !v_RM_5718_out0) || (!v_RD_3027_out0) && v_RM_5718_out0);
assign v_G2_6191_out0 = v_RD_3027_out0 && v_RM_5718_out0;
assign v_CARRY_2528_out0 = v_G2_6191_out0;
assign v_S_4515_out0 = v_G1_3946_out0;
assign v_S_671_out0 = v_S_4515_out0;
assign v_G1_2023_out0 = v_CARRY_2528_out0 || v_CARRY_2527_out0;
assign v_COUT_407_out0 = v_G1_2023_out0;
assign v__1369_out0 = { v__993_out0,v_S_671_out0 };
assign v_CIN_4912_out0 = v_COUT_407_out0;
assign v_RD_3037_out0 = v_CIN_4912_out0;
assign v_G1_3956_out0 = ((v_RD_3037_out0 && !v_RM_5728_out0) || (!v_RD_3037_out0) && v_RM_5728_out0);
assign v_G2_6201_out0 = v_RD_3037_out0 && v_RM_5728_out0;
assign v_CARRY_2538_out0 = v_G2_6201_out0;
assign v_S_4525_out0 = v_G1_3956_out0;
assign v_S_676_out0 = v_S_4525_out0;
assign v_G1_2028_out0 = v_CARRY_2538_out0 || v_CARRY_2537_out0;
assign v_COUT_412_out0 = v_G1_2028_out0;
assign v__896_out0 = { v__1369_out0,v_S_676_out0 };
assign v_CIN_4908_out0 = v_COUT_412_out0;
assign v_RD_3029_out0 = v_CIN_4908_out0;
assign v_G1_3948_out0 = ((v_RD_3029_out0 && !v_RM_5720_out0) || (!v_RD_3029_out0) && v_RM_5720_out0);
assign v_G2_6193_out0 = v_RD_3029_out0 && v_RM_5720_out0;
assign v_CARRY_2530_out0 = v_G2_6193_out0;
assign v_S_4517_out0 = v_G1_3948_out0;
assign v_S_672_out0 = v_S_4517_out0;
assign v_G1_2024_out0 = v_CARRY_2530_out0 || v_CARRY_2529_out0;
assign v_COUT_408_out0 = v_G1_2024_out0;
assign v__2225_out0 = { v__896_out0,v_S_672_out0 };
assign v_RM_1706_out0 = v_COUT_408_out0;
assign v_RM_5721_out0 = v_RM_1706_out0;
assign v_G1_3949_out0 = ((v_RD_3030_out0 && !v_RM_5721_out0) || (!v_RD_3030_out0) && v_RM_5721_out0);
assign v_G2_6194_out0 = v_RD_3030_out0 && v_RM_5721_out0;
assign v_CARRY_2531_out0 = v_G2_6194_out0;
assign v_S_4518_out0 = v_G1_3949_out0;
assign v_RM_5722_out0 = v_S_4518_out0;
assign v_G1_3950_out0 = ((v_RD_3031_out0 && !v_RM_5722_out0) || (!v_RD_3031_out0) && v_RM_5722_out0);
assign v_G2_6195_out0 = v_RD_3031_out0 && v_RM_5722_out0;
assign v_CARRY_2532_out0 = v_G2_6195_out0;
assign v_S_4519_out0 = v_G1_3950_out0;
assign v_S_673_out0 = v_S_4519_out0;
assign v_G1_2025_out0 = v_CARRY_2532_out0 || v_CARRY_2531_out0;
assign v_COUT_409_out0 = v_G1_2025_out0;
assign v__5248_out0 = { v__2225_out0,v_S_673_out0 };
assign v__5391_out0 = { v__5248_out0,v_COUT_409_out0 };
assign v_COUT_5376_out0 = v__5391_out0;
assign v_CIN_1150_out0 = v_COUT_5376_out0;
assign v__232_out0 = v_CIN_1150_out0[8:8];
assign v__870_out0 = v_CIN_1150_out0[6:6];
assign v__1053_out0 = v_CIN_1150_out0[3:3];
assign v__1072_out0 = v_CIN_1150_out0[15:15];
assign v__1223_out0 = v_CIN_1150_out0[0:0];
assign v__1491_out0 = v_CIN_1150_out0[9:9];
assign v__1507_out0 = v_CIN_1150_out0[2:2];
assign v__1533_out0 = v_CIN_1150_out0[7:7];
assign v__1866_out0 = v_CIN_1150_out0[1:1];
assign v__1884_out0 = v_CIN_1150_out0[10:10];
assign v__3343_out0 = v_CIN_1150_out0[11:11];
assign v__3759_out0 = v_CIN_1150_out0[12:12];
assign v__4285_out0 = v_CIN_1150_out0[13:13];
assign v__4318_out0 = v_CIN_1150_out0[14:14];
assign v__5279_out0 = v_CIN_1150_out0[5:5];
assign v__6627_out0 = v_CIN_1150_out0[4:4];
assign v_RM_1674_out0 = v__3759_out0;
assign v_RM_1675_out0 = v__4318_out0;
assign v_RM_1677_out0 = v__5279_out0;
assign v_RM_1678_out0 = v__6627_out0;
assign v_RM_1679_out0 = v__4285_out0;
assign v_RM_1680_out0 = v__1491_out0;
assign v_RM_1681_out0 = v__1884_out0;
assign v_RM_1682_out0 = v__1866_out0;
assign v_RM_1683_out0 = v__1053_out0;
assign v_RM_1684_out0 = v__870_out0;
assign v_RM_1685_out0 = v__1533_out0;
assign v_RM_1686_out0 = v__3343_out0;
assign v_RM_1687_out0 = v__232_out0;
assign v_RM_1688_out0 = v__1507_out0;
assign v_CIN_4879_out0 = v__1072_out0;
assign v_RM_5667_out0 = v__1223_out0;
assign v_RD_2969_out0 = v_CIN_4879_out0;
assign v_G1_3895_out0 = ((v_RD_2976_out0 && !v_RM_5667_out0) || (!v_RD_2976_out0) && v_RM_5667_out0);
assign v_RM_5655_out0 = v_RM_1674_out0;
assign v_RM_5657_out0 = v_RM_1675_out0;
assign v_RM_5661_out0 = v_RM_1677_out0;
assign v_RM_5663_out0 = v_RM_1678_out0;
assign v_RM_5665_out0 = v_RM_1679_out0;
assign v_RM_5668_out0 = v_RM_1680_out0;
assign v_RM_5670_out0 = v_RM_1681_out0;
assign v_RM_5672_out0 = v_RM_1682_out0;
assign v_RM_5674_out0 = v_RM_1683_out0;
assign v_RM_5676_out0 = v_RM_1684_out0;
assign v_RM_5678_out0 = v_RM_1685_out0;
assign v_RM_5680_out0 = v_RM_1686_out0;
assign v_RM_5682_out0 = v_RM_1687_out0;
assign v_RM_5684_out0 = v_RM_1688_out0;
assign v_G2_6140_out0 = v_RD_2976_out0 && v_RM_5667_out0;
assign v_CARRY_2477_out0 = v_G2_6140_out0;
assign v_G1_3883_out0 = ((v_RD_2964_out0 && !v_RM_5655_out0) || (!v_RD_2964_out0) && v_RM_5655_out0);
assign v_G1_3885_out0 = ((v_RD_2966_out0 && !v_RM_5657_out0) || (!v_RD_2966_out0) && v_RM_5657_out0);
assign v_G1_3889_out0 = ((v_RD_2970_out0 && !v_RM_5661_out0) || (!v_RD_2970_out0) && v_RM_5661_out0);
assign v_G1_3891_out0 = ((v_RD_2972_out0 && !v_RM_5663_out0) || (!v_RD_2972_out0) && v_RM_5663_out0);
assign v_G1_3893_out0 = ((v_RD_2974_out0 && !v_RM_5665_out0) || (!v_RD_2974_out0) && v_RM_5665_out0);
assign v_G1_3896_out0 = ((v_RD_2977_out0 && !v_RM_5668_out0) || (!v_RD_2977_out0) && v_RM_5668_out0);
assign v_G1_3898_out0 = ((v_RD_2979_out0 && !v_RM_5670_out0) || (!v_RD_2979_out0) && v_RM_5670_out0);
assign v_G1_3900_out0 = ((v_RD_2981_out0 && !v_RM_5672_out0) || (!v_RD_2981_out0) && v_RM_5672_out0);
assign v_G1_3902_out0 = ((v_RD_2983_out0 && !v_RM_5674_out0) || (!v_RD_2983_out0) && v_RM_5674_out0);
assign v_G1_3904_out0 = ((v_RD_2985_out0 && !v_RM_5676_out0) || (!v_RD_2985_out0) && v_RM_5676_out0);
assign v_G1_3906_out0 = ((v_RD_2987_out0 && !v_RM_5678_out0) || (!v_RD_2987_out0) && v_RM_5678_out0);
assign v_G1_3908_out0 = ((v_RD_2989_out0 && !v_RM_5680_out0) || (!v_RD_2989_out0) && v_RM_5680_out0);
assign v_G1_3910_out0 = ((v_RD_2991_out0 && !v_RM_5682_out0) || (!v_RD_2991_out0) && v_RM_5682_out0);
assign v_G1_3912_out0 = ((v_RD_2993_out0 && !v_RM_5684_out0) || (!v_RD_2993_out0) && v_RM_5684_out0);
assign v_S_4464_out0 = v_G1_3895_out0;
assign v_G2_6128_out0 = v_RD_2964_out0 && v_RM_5655_out0;
assign v_G2_6130_out0 = v_RD_2966_out0 && v_RM_5657_out0;
assign v_G2_6134_out0 = v_RD_2970_out0 && v_RM_5661_out0;
assign v_G2_6136_out0 = v_RD_2972_out0 && v_RM_5663_out0;
assign v_G2_6138_out0 = v_RD_2974_out0 && v_RM_5665_out0;
assign v_G2_6141_out0 = v_RD_2977_out0 && v_RM_5668_out0;
assign v_G2_6143_out0 = v_RD_2979_out0 && v_RM_5670_out0;
assign v_G2_6145_out0 = v_RD_2981_out0 && v_RM_5672_out0;
assign v_G2_6147_out0 = v_RD_2983_out0 && v_RM_5674_out0;
assign v_G2_6149_out0 = v_RD_2985_out0 && v_RM_5676_out0;
assign v_G2_6151_out0 = v_RD_2987_out0 && v_RM_5678_out0;
assign v_G2_6153_out0 = v_RD_2989_out0 && v_RM_5680_out0;
assign v_G2_6155_out0 = v_RD_2991_out0 && v_RM_5682_out0;
assign v_G2_6157_out0 = v_RD_2993_out0 && v_RM_5684_out0;
assign v_S_2281_out0 = v_S_4464_out0;
assign v_CARRY_2465_out0 = v_G2_6128_out0;
assign v_CARRY_2467_out0 = v_G2_6130_out0;
assign v_CARRY_2471_out0 = v_G2_6134_out0;
assign v_CARRY_2473_out0 = v_G2_6136_out0;
assign v_CARRY_2475_out0 = v_G2_6138_out0;
assign v_CARRY_2478_out0 = v_G2_6141_out0;
assign v_CARRY_2480_out0 = v_G2_6143_out0;
assign v_CARRY_2482_out0 = v_G2_6145_out0;
assign v_CARRY_2484_out0 = v_G2_6147_out0;
assign v_CARRY_2486_out0 = v_G2_6149_out0;
assign v_CARRY_2488_out0 = v_G2_6151_out0;
assign v_CARRY_2490_out0 = v_G2_6153_out0;
assign v_CARRY_2492_out0 = v_G2_6155_out0;
assign v_CARRY_2494_out0 = v_G2_6157_out0;
assign v_S_4452_out0 = v_G1_3883_out0;
assign v_S_4454_out0 = v_G1_3885_out0;
assign v_S_4458_out0 = v_G1_3889_out0;
assign v_S_4460_out0 = v_G1_3891_out0;
assign v_S_4462_out0 = v_G1_3893_out0;
assign v_S_4465_out0 = v_G1_3896_out0;
assign v_S_4467_out0 = v_G1_3898_out0;
assign v_S_4469_out0 = v_G1_3900_out0;
assign v_S_4471_out0 = v_G1_3902_out0;
assign v_S_4473_out0 = v_G1_3904_out0;
assign v_S_4475_out0 = v_G1_3906_out0;
assign v_S_4477_out0 = v_G1_3908_out0;
assign v_S_4479_out0 = v_G1_3910_out0;
assign v_S_4481_out0 = v_G1_3912_out0;
assign v_CIN_4885_out0 = v_CARRY_2477_out0;
assign v__1187_out0 = { v__1068_out0,v_S_2281_out0 };
assign v_RD_2982_out0 = v_CIN_4885_out0;
assign v_RM_5656_out0 = v_S_4452_out0;
assign v_RM_5658_out0 = v_S_4454_out0;
assign v_RM_5662_out0 = v_S_4458_out0;
assign v_RM_5664_out0 = v_S_4460_out0;
assign v_RM_5666_out0 = v_S_4462_out0;
assign v_RM_5669_out0 = v_S_4465_out0;
assign v_RM_5671_out0 = v_S_4467_out0;
assign v_RM_5673_out0 = v_S_4469_out0;
assign v_RM_5675_out0 = v_S_4471_out0;
assign v_RM_5677_out0 = v_S_4473_out0;
assign v_RM_5679_out0 = v_S_4475_out0;
assign v_RM_5681_out0 = v_S_4477_out0;
assign v_RM_5683_out0 = v_S_4479_out0;
assign v_RM_5685_out0 = v_S_4481_out0;
assign v_G1_3901_out0 = ((v_RD_2982_out0 && !v_RM_5673_out0) || (!v_RD_2982_out0) && v_RM_5673_out0);
assign v_G2_6146_out0 = v_RD_2982_out0 && v_RM_5673_out0;
assign v_CARRY_2483_out0 = v_G2_6146_out0;
assign v_S_4470_out0 = v_G1_3901_out0;
assign v_S_649_out0 = v_S_4470_out0;
assign v_G1_2001_out0 = v_CARRY_2483_out0 || v_CARRY_2482_out0;
assign v_COUT_385_out0 = v_G1_2001_out0;
assign v_CIN_4891_out0 = v_COUT_385_out0;
assign v_RD_2994_out0 = v_CIN_4891_out0;
assign v_G1_3913_out0 = ((v_RD_2994_out0 && !v_RM_5685_out0) || (!v_RD_2994_out0) && v_RM_5685_out0);
assign v_G2_6158_out0 = v_RD_2994_out0 && v_RM_5685_out0;
assign v_CARRY_2495_out0 = v_G2_6158_out0;
assign v_S_4482_out0 = v_G1_3913_out0;
assign v_S_655_out0 = v_S_4482_out0;
assign v_G1_2007_out0 = v_CARRY_2495_out0 || v_CARRY_2494_out0;
assign v_COUT_391_out0 = v_G1_2007_out0;
assign v__2338_out0 = { v_S_649_out0,v_S_655_out0 };
assign v_CIN_4886_out0 = v_COUT_391_out0;
assign v_RD_2984_out0 = v_CIN_4886_out0;
assign v_G1_3903_out0 = ((v_RD_2984_out0 && !v_RM_5675_out0) || (!v_RD_2984_out0) && v_RM_5675_out0);
assign v_G2_6148_out0 = v_RD_2984_out0 && v_RM_5675_out0;
assign v_CARRY_2485_out0 = v_G2_6148_out0;
assign v_S_4472_out0 = v_G1_3903_out0;
assign v_S_650_out0 = v_S_4472_out0;
assign v_G1_2002_out0 = v_CARRY_2485_out0 || v_CARRY_2484_out0;
assign v_COUT_386_out0 = v_G1_2002_out0;
assign v__1247_out0 = { v__2338_out0,v_S_650_out0 };
assign v_CIN_4881_out0 = v_COUT_386_out0;
assign v_RD_2973_out0 = v_CIN_4881_out0;
assign v_G1_3892_out0 = ((v_RD_2973_out0 && !v_RM_5664_out0) || (!v_RD_2973_out0) && v_RM_5664_out0);
assign v_G2_6137_out0 = v_RD_2973_out0 && v_RM_5664_out0;
assign v_CARRY_2474_out0 = v_G2_6137_out0;
assign v_S_4461_out0 = v_G1_3892_out0;
assign v_S_645_out0 = v_S_4461_out0;
assign v_G1_1997_out0 = v_CARRY_2474_out0 || v_CARRY_2473_out0;
assign v_COUT_381_out0 = v_G1_1997_out0;
assign v__3455_out0 = { v__1247_out0,v_S_645_out0 };
assign v_CIN_4880_out0 = v_COUT_381_out0;
assign v_RD_2971_out0 = v_CIN_4880_out0;
assign v_G1_3890_out0 = ((v_RD_2971_out0 && !v_RM_5662_out0) || (!v_RD_2971_out0) && v_RM_5662_out0);
assign v_G2_6135_out0 = v_RD_2971_out0 && v_RM_5662_out0;
assign v_CARRY_2472_out0 = v_G2_6135_out0;
assign v_S_4459_out0 = v_G1_3890_out0;
assign v_S_644_out0 = v_S_4459_out0;
assign v_G1_1996_out0 = v_CARRY_2472_out0 || v_CARRY_2471_out0;
assign v_COUT_380_out0 = v_G1_1996_out0;
assign v__6665_out0 = { v__3455_out0,v_S_644_out0 };
assign v_CIN_4887_out0 = v_COUT_380_out0;
assign v_RD_2986_out0 = v_CIN_4887_out0;
assign v_G1_3905_out0 = ((v_RD_2986_out0 && !v_RM_5677_out0) || (!v_RD_2986_out0) && v_RM_5677_out0);
assign v_G2_6150_out0 = v_RD_2986_out0 && v_RM_5677_out0;
assign v_CARRY_2487_out0 = v_G2_6150_out0;
assign v_S_4474_out0 = v_G1_3905_out0;
assign v_S_651_out0 = v_S_4474_out0;
assign v_G1_2003_out0 = v_CARRY_2487_out0 || v_CARRY_2486_out0;
assign v_COUT_387_out0 = v_G1_2003_out0;
assign v__1613_out0 = { v__6665_out0,v_S_651_out0 };
assign v_CIN_4888_out0 = v_COUT_387_out0;
assign v_RD_2988_out0 = v_CIN_4888_out0;
assign v_G1_3907_out0 = ((v_RD_2988_out0 && !v_RM_5679_out0) || (!v_RD_2988_out0) && v_RM_5679_out0);
assign v_G2_6152_out0 = v_RD_2988_out0 && v_RM_5679_out0;
assign v_CARRY_2489_out0 = v_G2_6152_out0;
assign v_S_4476_out0 = v_G1_3907_out0;
assign v_S_652_out0 = v_S_4476_out0;
assign v_G1_2004_out0 = v_CARRY_2489_out0 || v_CARRY_2488_out0;
assign v_COUT_388_out0 = v_G1_2004_out0;
assign v__3510_out0 = { v__1613_out0,v_S_652_out0 };
assign v_CIN_4890_out0 = v_COUT_388_out0;
assign v_RD_2992_out0 = v_CIN_4890_out0;
assign v_G1_3911_out0 = ((v_RD_2992_out0 && !v_RM_5683_out0) || (!v_RD_2992_out0) && v_RM_5683_out0);
assign v_G2_6156_out0 = v_RD_2992_out0 && v_RM_5683_out0;
assign v_CARRY_2493_out0 = v_G2_6156_out0;
assign v_S_4480_out0 = v_G1_3911_out0;
assign v_S_654_out0 = v_S_4480_out0;
assign v_G1_2006_out0 = v_CARRY_2493_out0 || v_CARRY_2492_out0;
assign v_COUT_390_out0 = v_G1_2006_out0;
assign v__2321_out0 = { v__3510_out0,v_S_654_out0 };
assign v_CIN_4883_out0 = v_COUT_390_out0;
assign v_RD_2978_out0 = v_CIN_4883_out0;
assign v_G1_3897_out0 = ((v_RD_2978_out0 && !v_RM_5669_out0) || (!v_RD_2978_out0) && v_RM_5669_out0);
assign v_G2_6142_out0 = v_RD_2978_out0 && v_RM_5669_out0;
assign v_CARRY_2479_out0 = v_G2_6142_out0;
assign v_S_4466_out0 = v_G1_3897_out0;
assign v_S_647_out0 = v_S_4466_out0;
assign v_G1_1999_out0 = v_CARRY_2479_out0 || v_CARRY_2478_out0;
assign v_COUT_383_out0 = v_G1_1999_out0;
assign v__3403_out0 = { v__2321_out0,v_S_647_out0 };
assign v_CIN_4884_out0 = v_COUT_383_out0;
assign v_RD_2980_out0 = v_CIN_4884_out0;
assign v_G1_3899_out0 = ((v_RD_2980_out0 && !v_RM_5671_out0) || (!v_RD_2980_out0) && v_RM_5671_out0);
assign v_G2_6144_out0 = v_RD_2980_out0 && v_RM_5671_out0;
assign v_CARRY_2481_out0 = v_G2_6144_out0;
assign v_S_4468_out0 = v_G1_3899_out0;
assign v_S_648_out0 = v_S_4468_out0;
assign v_G1_2000_out0 = v_CARRY_2481_out0 || v_CARRY_2480_out0;
assign v_COUT_384_out0 = v_G1_2000_out0;
assign v__2847_out0 = { v__3403_out0,v_S_648_out0 };
assign v_CIN_4889_out0 = v_COUT_384_out0;
assign v_RD_2990_out0 = v_CIN_4889_out0;
assign v_G1_3909_out0 = ((v_RD_2990_out0 && !v_RM_5681_out0) || (!v_RD_2990_out0) && v_RM_5681_out0);
assign v_G2_6154_out0 = v_RD_2990_out0 && v_RM_5681_out0;
assign v_CARRY_2491_out0 = v_G2_6154_out0;
assign v_S_4478_out0 = v_G1_3909_out0;
assign v_S_653_out0 = v_S_4478_out0;
assign v_G1_2005_out0 = v_CARRY_2491_out0 || v_CARRY_2490_out0;
assign v_COUT_389_out0 = v_G1_2005_out0;
assign v__991_out0 = { v__2847_out0,v_S_653_out0 };
assign v_CIN_4877_out0 = v_COUT_389_out0;
assign v_RD_2965_out0 = v_CIN_4877_out0;
assign v_G1_3884_out0 = ((v_RD_2965_out0 && !v_RM_5656_out0) || (!v_RD_2965_out0) && v_RM_5656_out0);
assign v_G2_6129_out0 = v_RD_2965_out0 && v_RM_5656_out0;
assign v_CARRY_2466_out0 = v_G2_6129_out0;
assign v_S_4453_out0 = v_G1_3884_out0;
assign v_S_641_out0 = v_S_4453_out0;
assign v_G1_1993_out0 = v_CARRY_2466_out0 || v_CARRY_2465_out0;
assign v_COUT_377_out0 = v_G1_1993_out0;
assign v__1367_out0 = { v__991_out0,v_S_641_out0 };
assign v_CIN_4882_out0 = v_COUT_377_out0;
assign v_RD_2975_out0 = v_CIN_4882_out0;
assign v_G1_3894_out0 = ((v_RD_2975_out0 && !v_RM_5666_out0) || (!v_RD_2975_out0) && v_RM_5666_out0);
assign v_G2_6139_out0 = v_RD_2975_out0 && v_RM_5666_out0;
assign v_CARRY_2476_out0 = v_G2_6139_out0;
assign v_S_4463_out0 = v_G1_3894_out0;
assign v_S_646_out0 = v_S_4463_out0;
assign v_G1_1998_out0 = v_CARRY_2476_out0 || v_CARRY_2475_out0;
assign v_COUT_382_out0 = v_G1_1998_out0;
assign v__894_out0 = { v__1367_out0,v_S_646_out0 };
assign v_CIN_4878_out0 = v_COUT_382_out0;
assign v_RD_2967_out0 = v_CIN_4878_out0;
assign v_G1_3886_out0 = ((v_RD_2967_out0 && !v_RM_5658_out0) || (!v_RD_2967_out0) && v_RM_5658_out0);
assign v_G2_6131_out0 = v_RD_2967_out0 && v_RM_5658_out0;
assign v_CARRY_2468_out0 = v_G2_6131_out0;
assign v_S_4455_out0 = v_G1_3886_out0;
assign v_S_642_out0 = v_S_4455_out0;
assign v_G1_1994_out0 = v_CARRY_2468_out0 || v_CARRY_2467_out0;
assign v_COUT_378_out0 = v_G1_1994_out0;
assign v__2223_out0 = { v__894_out0,v_S_642_out0 };
assign v_RM_1676_out0 = v_COUT_378_out0;
assign v_RM_5659_out0 = v_RM_1676_out0;
assign v_G1_3887_out0 = ((v_RD_2968_out0 && !v_RM_5659_out0) || (!v_RD_2968_out0) && v_RM_5659_out0);
assign v_G2_6132_out0 = v_RD_2968_out0 && v_RM_5659_out0;
assign v_CARRY_2469_out0 = v_G2_6132_out0;
assign v_S_4456_out0 = v_G1_3887_out0;
assign v_RM_5660_out0 = v_S_4456_out0;
assign v_G1_3888_out0 = ((v_RD_2969_out0 && !v_RM_5660_out0) || (!v_RD_2969_out0) && v_RM_5660_out0);
assign v_G2_6133_out0 = v_RD_2969_out0 && v_RM_5660_out0;
assign v_CARRY_2470_out0 = v_G2_6133_out0;
assign v_S_4457_out0 = v_G1_3888_out0;
assign v_S_643_out0 = v_S_4457_out0;
assign v_G1_1995_out0 = v_CARRY_2470_out0 || v_CARRY_2469_out0;
assign v_COUT_379_out0 = v_G1_1995_out0;
assign v__5246_out0 = { v__2223_out0,v_S_643_out0 };
assign v__5389_out0 = { v__5246_out0,v_COUT_379_out0 };
assign v_COUT_5374_out0 = v__5389_out0;
assign v_CIN_1155_out0 = v_COUT_5374_out0;
assign v__237_out0 = v_CIN_1155_out0[8:8];
assign v__875_out0 = v_CIN_1155_out0[6:6];
assign v__1058_out0 = v_CIN_1155_out0[3:3];
assign v__1077_out0 = v_CIN_1155_out0[15:15];
assign v__1228_out0 = v_CIN_1155_out0[0:0];
assign v__1496_out0 = v_CIN_1155_out0[9:9];
assign v__1512_out0 = v_CIN_1155_out0[2:2];
assign v__1538_out0 = v_CIN_1155_out0[7:7];
assign v__1871_out0 = v_CIN_1155_out0[1:1];
assign v__1889_out0 = v_CIN_1155_out0[10:10];
assign v__3348_out0 = v_CIN_1155_out0[11:11];
assign v__3764_out0 = v_CIN_1155_out0[12:12];
assign v__4290_out0 = v_CIN_1155_out0[13:13];
assign v__4323_out0 = v_CIN_1155_out0[14:14];
assign v__5284_out0 = v_CIN_1155_out0[5:5];
assign v__6632_out0 = v_CIN_1155_out0[4:4];
assign v_RM_1749_out0 = v__3764_out0;
assign v_RM_1750_out0 = v__4323_out0;
assign v_RM_1752_out0 = v__5284_out0;
assign v_RM_1753_out0 = v__6632_out0;
assign v_RM_1754_out0 = v__4290_out0;
assign v_RM_1755_out0 = v__1496_out0;
assign v_RM_1756_out0 = v__1889_out0;
assign v_RM_1757_out0 = v__1871_out0;
assign v_RM_1758_out0 = v__1058_out0;
assign v_RM_1759_out0 = v__875_out0;
assign v_RM_1760_out0 = v__1538_out0;
assign v_RM_1761_out0 = v__3348_out0;
assign v_RM_1762_out0 = v__237_out0;
assign v_RM_1763_out0 = v__1512_out0;
assign v_CIN_4954_out0 = v__1077_out0;
assign v_RM_5822_out0 = v__1228_out0;
assign v_RD_3124_out0 = v_CIN_4954_out0;
assign v_G1_4050_out0 = ((v_RD_3131_out0 && !v_RM_5822_out0) || (!v_RD_3131_out0) && v_RM_5822_out0);
assign v_RM_5810_out0 = v_RM_1749_out0;
assign v_RM_5812_out0 = v_RM_1750_out0;
assign v_RM_5816_out0 = v_RM_1752_out0;
assign v_RM_5818_out0 = v_RM_1753_out0;
assign v_RM_5820_out0 = v_RM_1754_out0;
assign v_RM_5823_out0 = v_RM_1755_out0;
assign v_RM_5825_out0 = v_RM_1756_out0;
assign v_RM_5827_out0 = v_RM_1757_out0;
assign v_RM_5829_out0 = v_RM_1758_out0;
assign v_RM_5831_out0 = v_RM_1759_out0;
assign v_RM_5833_out0 = v_RM_1760_out0;
assign v_RM_5835_out0 = v_RM_1761_out0;
assign v_RM_5837_out0 = v_RM_1762_out0;
assign v_RM_5839_out0 = v_RM_1763_out0;
assign v_G2_6295_out0 = v_RD_3131_out0 && v_RM_5822_out0;
assign v_CARRY_2632_out0 = v_G2_6295_out0;
assign v_G1_4038_out0 = ((v_RD_3119_out0 && !v_RM_5810_out0) || (!v_RD_3119_out0) && v_RM_5810_out0);
assign v_G1_4040_out0 = ((v_RD_3121_out0 && !v_RM_5812_out0) || (!v_RD_3121_out0) && v_RM_5812_out0);
assign v_G1_4044_out0 = ((v_RD_3125_out0 && !v_RM_5816_out0) || (!v_RD_3125_out0) && v_RM_5816_out0);
assign v_G1_4046_out0 = ((v_RD_3127_out0 && !v_RM_5818_out0) || (!v_RD_3127_out0) && v_RM_5818_out0);
assign v_G1_4048_out0 = ((v_RD_3129_out0 && !v_RM_5820_out0) || (!v_RD_3129_out0) && v_RM_5820_out0);
assign v_G1_4051_out0 = ((v_RD_3132_out0 && !v_RM_5823_out0) || (!v_RD_3132_out0) && v_RM_5823_out0);
assign v_G1_4053_out0 = ((v_RD_3134_out0 && !v_RM_5825_out0) || (!v_RD_3134_out0) && v_RM_5825_out0);
assign v_G1_4055_out0 = ((v_RD_3136_out0 && !v_RM_5827_out0) || (!v_RD_3136_out0) && v_RM_5827_out0);
assign v_G1_4057_out0 = ((v_RD_3138_out0 && !v_RM_5829_out0) || (!v_RD_3138_out0) && v_RM_5829_out0);
assign v_G1_4059_out0 = ((v_RD_3140_out0 && !v_RM_5831_out0) || (!v_RD_3140_out0) && v_RM_5831_out0);
assign v_G1_4061_out0 = ((v_RD_3142_out0 && !v_RM_5833_out0) || (!v_RD_3142_out0) && v_RM_5833_out0);
assign v_G1_4063_out0 = ((v_RD_3144_out0 && !v_RM_5835_out0) || (!v_RD_3144_out0) && v_RM_5835_out0);
assign v_G1_4065_out0 = ((v_RD_3146_out0 && !v_RM_5837_out0) || (!v_RD_3146_out0) && v_RM_5837_out0);
assign v_G1_4067_out0 = ((v_RD_3148_out0 && !v_RM_5839_out0) || (!v_RD_3148_out0) && v_RM_5839_out0);
assign v_S_4619_out0 = v_G1_4050_out0;
assign v_G2_6283_out0 = v_RD_3119_out0 && v_RM_5810_out0;
assign v_G2_6285_out0 = v_RD_3121_out0 && v_RM_5812_out0;
assign v_G2_6289_out0 = v_RD_3125_out0 && v_RM_5816_out0;
assign v_G2_6291_out0 = v_RD_3127_out0 && v_RM_5818_out0;
assign v_G2_6293_out0 = v_RD_3129_out0 && v_RM_5820_out0;
assign v_G2_6296_out0 = v_RD_3132_out0 && v_RM_5823_out0;
assign v_G2_6298_out0 = v_RD_3134_out0 && v_RM_5825_out0;
assign v_G2_6300_out0 = v_RD_3136_out0 && v_RM_5827_out0;
assign v_G2_6302_out0 = v_RD_3138_out0 && v_RM_5829_out0;
assign v_G2_6304_out0 = v_RD_3140_out0 && v_RM_5831_out0;
assign v_G2_6306_out0 = v_RD_3142_out0 && v_RM_5833_out0;
assign v_G2_6308_out0 = v_RD_3144_out0 && v_RM_5835_out0;
assign v_G2_6310_out0 = v_RD_3146_out0 && v_RM_5837_out0;
assign v_G2_6312_out0 = v_RD_3148_out0 && v_RM_5839_out0;
assign v_S_2286_out0 = v_S_4619_out0;
assign v_CARRY_2620_out0 = v_G2_6283_out0;
assign v_CARRY_2622_out0 = v_G2_6285_out0;
assign v_CARRY_2626_out0 = v_G2_6289_out0;
assign v_CARRY_2628_out0 = v_G2_6291_out0;
assign v_CARRY_2630_out0 = v_G2_6293_out0;
assign v_CARRY_2633_out0 = v_G2_6296_out0;
assign v_CARRY_2635_out0 = v_G2_6298_out0;
assign v_CARRY_2637_out0 = v_G2_6300_out0;
assign v_CARRY_2639_out0 = v_G2_6302_out0;
assign v_CARRY_2641_out0 = v_G2_6304_out0;
assign v_CARRY_2643_out0 = v_G2_6306_out0;
assign v_CARRY_2645_out0 = v_G2_6308_out0;
assign v_CARRY_2647_out0 = v_G2_6310_out0;
assign v_CARRY_2649_out0 = v_G2_6312_out0;
assign v_S_4607_out0 = v_G1_4038_out0;
assign v_S_4609_out0 = v_G1_4040_out0;
assign v_S_4613_out0 = v_G1_4044_out0;
assign v_S_4615_out0 = v_G1_4046_out0;
assign v_S_4617_out0 = v_G1_4048_out0;
assign v_S_4620_out0 = v_G1_4051_out0;
assign v_S_4622_out0 = v_G1_4053_out0;
assign v_S_4624_out0 = v_G1_4055_out0;
assign v_S_4626_out0 = v_G1_4057_out0;
assign v_S_4628_out0 = v_G1_4059_out0;
assign v_S_4630_out0 = v_G1_4061_out0;
assign v_S_4632_out0 = v_G1_4063_out0;
assign v_S_4634_out0 = v_G1_4065_out0;
assign v_S_4636_out0 = v_G1_4067_out0;
assign v_CIN_4960_out0 = v_CARRY_2632_out0;
assign v_RD_3137_out0 = v_CIN_4960_out0;
assign v__4830_out0 = { v__1187_out0,v_S_2286_out0 };
assign v_RM_5811_out0 = v_S_4607_out0;
assign v_RM_5813_out0 = v_S_4609_out0;
assign v_RM_5817_out0 = v_S_4613_out0;
assign v_RM_5819_out0 = v_S_4615_out0;
assign v_RM_5821_out0 = v_S_4617_out0;
assign v_RM_5824_out0 = v_S_4620_out0;
assign v_RM_5826_out0 = v_S_4622_out0;
assign v_RM_5828_out0 = v_S_4624_out0;
assign v_RM_5830_out0 = v_S_4626_out0;
assign v_RM_5832_out0 = v_S_4628_out0;
assign v_RM_5834_out0 = v_S_4630_out0;
assign v_RM_5836_out0 = v_S_4632_out0;
assign v_RM_5838_out0 = v_S_4634_out0;
assign v_RM_5840_out0 = v_S_4636_out0;
assign v_G1_4056_out0 = ((v_RD_3137_out0 && !v_RM_5828_out0) || (!v_RD_3137_out0) && v_RM_5828_out0);
assign v_G2_6301_out0 = v_RD_3137_out0 && v_RM_5828_out0;
assign v_CARRY_2638_out0 = v_G2_6301_out0;
assign v_S_4625_out0 = v_G1_4056_out0;
assign v_S_724_out0 = v_S_4625_out0;
assign v_G1_2076_out0 = v_CARRY_2638_out0 || v_CARRY_2637_out0;
assign v_COUT_460_out0 = v_G1_2076_out0;
assign v_CIN_4966_out0 = v_COUT_460_out0;
assign v_RD_3149_out0 = v_CIN_4966_out0;
assign v_G1_4068_out0 = ((v_RD_3149_out0 && !v_RM_5840_out0) || (!v_RD_3149_out0) && v_RM_5840_out0);
assign v_G2_6313_out0 = v_RD_3149_out0 && v_RM_5840_out0;
assign v_CARRY_2650_out0 = v_G2_6313_out0;
assign v_S_4637_out0 = v_G1_4068_out0;
assign v_S_730_out0 = v_S_4637_out0;
assign v_G1_2082_out0 = v_CARRY_2650_out0 || v_CARRY_2649_out0;
assign v_COUT_466_out0 = v_G1_2082_out0;
assign v__2343_out0 = { v_S_724_out0,v_S_730_out0 };
assign v_CIN_4961_out0 = v_COUT_466_out0;
assign v_RD_3139_out0 = v_CIN_4961_out0;
assign v_G1_4058_out0 = ((v_RD_3139_out0 && !v_RM_5830_out0) || (!v_RD_3139_out0) && v_RM_5830_out0);
assign v_G2_6303_out0 = v_RD_3139_out0 && v_RM_5830_out0;
assign v_CARRY_2640_out0 = v_G2_6303_out0;
assign v_S_4627_out0 = v_G1_4058_out0;
assign v_S_725_out0 = v_S_4627_out0;
assign v_G1_2077_out0 = v_CARRY_2640_out0 || v_CARRY_2639_out0;
assign v_COUT_461_out0 = v_G1_2077_out0;
assign v__1252_out0 = { v__2343_out0,v_S_725_out0 };
assign v_CIN_4956_out0 = v_COUT_461_out0;
assign v_RD_3128_out0 = v_CIN_4956_out0;
assign v_G1_4047_out0 = ((v_RD_3128_out0 && !v_RM_5819_out0) || (!v_RD_3128_out0) && v_RM_5819_out0);
assign v_G2_6292_out0 = v_RD_3128_out0 && v_RM_5819_out0;
assign v_CARRY_2629_out0 = v_G2_6292_out0;
assign v_S_4616_out0 = v_G1_4047_out0;
assign v_S_720_out0 = v_S_4616_out0;
assign v_G1_2072_out0 = v_CARRY_2629_out0 || v_CARRY_2628_out0;
assign v_COUT_456_out0 = v_G1_2072_out0;
assign v__3460_out0 = { v__1252_out0,v_S_720_out0 };
assign v_CIN_4955_out0 = v_COUT_456_out0;
assign v_RD_3126_out0 = v_CIN_4955_out0;
assign v_G1_4045_out0 = ((v_RD_3126_out0 && !v_RM_5817_out0) || (!v_RD_3126_out0) && v_RM_5817_out0);
assign v_G2_6290_out0 = v_RD_3126_out0 && v_RM_5817_out0;
assign v_CARRY_2627_out0 = v_G2_6290_out0;
assign v_S_4614_out0 = v_G1_4045_out0;
assign v_S_719_out0 = v_S_4614_out0;
assign v_G1_2071_out0 = v_CARRY_2627_out0 || v_CARRY_2626_out0;
assign v_COUT_455_out0 = v_G1_2071_out0;
assign v__6670_out0 = { v__3460_out0,v_S_719_out0 };
assign v_CIN_4962_out0 = v_COUT_455_out0;
assign v_RD_3141_out0 = v_CIN_4962_out0;
assign v_G1_4060_out0 = ((v_RD_3141_out0 && !v_RM_5832_out0) || (!v_RD_3141_out0) && v_RM_5832_out0);
assign v_G2_6305_out0 = v_RD_3141_out0 && v_RM_5832_out0;
assign v_CARRY_2642_out0 = v_G2_6305_out0;
assign v_S_4629_out0 = v_G1_4060_out0;
assign v_S_726_out0 = v_S_4629_out0;
assign v_G1_2078_out0 = v_CARRY_2642_out0 || v_CARRY_2641_out0;
assign v_COUT_462_out0 = v_G1_2078_out0;
assign v__1618_out0 = { v__6670_out0,v_S_726_out0 };
assign v_CIN_4963_out0 = v_COUT_462_out0;
assign v_RD_3143_out0 = v_CIN_4963_out0;
assign v_G1_4062_out0 = ((v_RD_3143_out0 && !v_RM_5834_out0) || (!v_RD_3143_out0) && v_RM_5834_out0);
assign v_G2_6307_out0 = v_RD_3143_out0 && v_RM_5834_out0;
assign v_CARRY_2644_out0 = v_G2_6307_out0;
assign v_S_4631_out0 = v_G1_4062_out0;
assign v_S_727_out0 = v_S_4631_out0;
assign v_G1_2079_out0 = v_CARRY_2644_out0 || v_CARRY_2643_out0;
assign v_COUT_463_out0 = v_G1_2079_out0;
assign v__3515_out0 = { v__1618_out0,v_S_727_out0 };
assign v_CIN_4965_out0 = v_COUT_463_out0;
assign v_RD_3147_out0 = v_CIN_4965_out0;
assign v_G1_4066_out0 = ((v_RD_3147_out0 && !v_RM_5838_out0) || (!v_RD_3147_out0) && v_RM_5838_out0);
assign v_G2_6311_out0 = v_RD_3147_out0 && v_RM_5838_out0;
assign v_CARRY_2648_out0 = v_G2_6311_out0;
assign v_S_4635_out0 = v_G1_4066_out0;
assign v_S_729_out0 = v_S_4635_out0;
assign v_G1_2081_out0 = v_CARRY_2648_out0 || v_CARRY_2647_out0;
assign v_COUT_465_out0 = v_G1_2081_out0;
assign v__2326_out0 = { v__3515_out0,v_S_729_out0 };
assign v_CIN_4958_out0 = v_COUT_465_out0;
assign v_RD_3133_out0 = v_CIN_4958_out0;
assign v_G1_4052_out0 = ((v_RD_3133_out0 && !v_RM_5824_out0) || (!v_RD_3133_out0) && v_RM_5824_out0);
assign v_G2_6297_out0 = v_RD_3133_out0 && v_RM_5824_out0;
assign v_CARRY_2634_out0 = v_G2_6297_out0;
assign v_S_4621_out0 = v_G1_4052_out0;
assign v_S_722_out0 = v_S_4621_out0;
assign v_G1_2074_out0 = v_CARRY_2634_out0 || v_CARRY_2633_out0;
assign v_COUT_458_out0 = v_G1_2074_out0;
assign v__3408_out0 = { v__2326_out0,v_S_722_out0 };
assign v_CIN_4959_out0 = v_COUT_458_out0;
assign v_RD_3135_out0 = v_CIN_4959_out0;
assign v_G1_4054_out0 = ((v_RD_3135_out0 && !v_RM_5826_out0) || (!v_RD_3135_out0) && v_RM_5826_out0);
assign v_G2_6299_out0 = v_RD_3135_out0 && v_RM_5826_out0;
assign v_CARRY_2636_out0 = v_G2_6299_out0;
assign v_S_4623_out0 = v_G1_4054_out0;
assign v_S_723_out0 = v_S_4623_out0;
assign v_G1_2075_out0 = v_CARRY_2636_out0 || v_CARRY_2635_out0;
assign v_COUT_459_out0 = v_G1_2075_out0;
assign v__2852_out0 = { v__3408_out0,v_S_723_out0 };
assign v_CIN_4964_out0 = v_COUT_459_out0;
assign v_RD_3145_out0 = v_CIN_4964_out0;
assign v_G1_4064_out0 = ((v_RD_3145_out0 && !v_RM_5836_out0) || (!v_RD_3145_out0) && v_RM_5836_out0);
assign v_G2_6309_out0 = v_RD_3145_out0 && v_RM_5836_out0;
assign v_CARRY_2646_out0 = v_G2_6309_out0;
assign v_S_4633_out0 = v_G1_4064_out0;
assign v_S_728_out0 = v_S_4633_out0;
assign v_G1_2080_out0 = v_CARRY_2646_out0 || v_CARRY_2645_out0;
assign v_COUT_464_out0 = v_G1_2080_out0;
assign v__996_out0 = { v__2852_out0,v_S_728_out0 };
assign v_CIN_4952_out0 = v_COUT_464_out0;
assign v_RD_3120_out0 = v_CIN_4952_out0;
assign v_G1_4039_out0 = ((v_RD_3120_out0 && !v_RM_5811_out0) || (!v_RD_3120_out0) && v_RM_5811_out0);
assign v_G2_6284_out0 = v_RD_3120_out0 && v_RM_5811_out0;
assign v_CARRY_2621_out0 = v_G2_6284_out0;
assign v_S_4608_out0 = v_G1_4039_out0;
assign v_S_716_out0 = v_S_4608_out0;
assign v_G1_2068_out0 = v_CARRY_2621_out0 || v_CARRY_2620_out0;
assign v_COUT_452_out0 = v_G1_2068_out0;
assign v__1372_out0 = { v__996_out0,v_S_716_out0 };
assign v_CIN_4957_out0 = v_COUT_452_out0;
assign v_RD_3130_out0 = v_CIN_4957_out0;
assign v_G1_4049_out0 = ((v_RD_3130_out0 && !v_RM_5821_out0) || (!v_RD_3130_out0) && v_RM_5821_out0);
assign v_G2_6294_out0 = v_RD_3130_out0 && v_RM_5821_out0;
assign v_CARRY_2631_out0 = v_G2_6294_out0;
assign v_S_4618_out0 = v_G1_4049_out0;
assign v_S_721_out0 = v_S_4618_out0;
assign v_G1_2073_out0 = v_CARRY_2631_out0 || v_CARRY_2630_out0;
assign v_COUT_457_out0 = v_G1_2073_out0;
assign v__899_out0 = { v__1372_out0,v_S_721_out0 };
assign v_CIN_4953_out0 = v_COUT_457_out0;
assign v_RD_3122_out0 = v_CIN_4953_out0;
assign v_G1_4041_out0 = ((v_RD_3122_out0 && !v_RM_5813_out0) || (!v_RD_3122_out0) && v_RM_5813_out0);
assign v_G2_6286_out0 = v_RD_3122_out0 && v_RM_5813_out0;
assign v_CARRY_2623_out0 = v_G2_6286_out0;
assign v_S_4610_out0 = v_G1_4041_out0;
assign v_S_717_out0 = v_S_4610_out0;
assign v_G1_2069_out0 = v_CARRY_2623_out0 || v_CARRY_2622_out0;
assign v_COUT_453_out0 = v_G1_2069_out0;
assign v__2228_out0 = { v__899_out0,v_S_717_out0 };
assign v_RM_1751_out0 = v_COUT_453_out0;
assign v_RM_5814_out0 = v_RM_1751_out0;
assign v_G1_4042_out0 = ((v_RD_3123_out0 && !v_RM_5814_out0) || (!v_RD_3123_out0) && v_RM_5814_out0);
assign v_G2_6287_out0 = v_RD_3123_out0 && v_RM_5814_out0;
assign v_CARRY_2624_out0 = v_G2_6287_out0;
assign v_S_4611_out0 = v_G1_4042_out0;
assign v_RM_5815_out0 = v_S_4611_out0;
assign v_G1_4043_out0 = ((v_RD_3124_out0 && !v_RM_5815_out0) || (!v_RD_3124_out0) && v_RM_5815_out0);
assign v_G2_6288_out0 = v_RD_3124_out0 && v_RM_5815_out0;
assign v_CARRY_2625_out0 = v_G2_6288_out0;
assign v_S_4612_out0 = v_G1_4043_out0;
assign v_S_718_out0 = v_S_4612_out0;
assign v_G1_2070_out0 = v_CARRY_2625_out0 || v_CARRY_2624_out0;
assign v_COUT_454_out0 = v_G1_2070_out0;
assign v__5251_out0 = { v__2228_out0,v_S_718_out0 };
assign v__5394_out0 = { v__5251_out0,v_COUT_454_out0 };
assign v_COUT_5379_out0 = v__5394_out0;
assign v_CIN_1159_out0 = v_COUT_5379_out0;
assign v__241_out0 = v_CIN_1159_out0[8:8];
assign v__879_out0 = v_CIN_1159_out0[6:6];
assign v__1062_out0 = v_CIN_1159_out0[3:3];
assign v__1081_out0 = v_CIN_1159_out0[15:15];
assign v__1232_out0 = v_CIN_1159_out0[0:0];
assign v__1500_out0 = v_CIN_1159_out0[9:9];
assign v__1516_out0 = v_CIN_1159_out0[2:2];
assign v__1542_out0 = v_CIN_1159_out0[7:7];
assign v__1875_out0 = v_CIN_1159_out0[1:1];
assign v__1893_out0 = v_CIN_1159_out0[10:10];
assign v__3352_out0 = v_CIN_1159_out0[11:11];
assign v__3768_out0 = v_CIN_1159_out0[12:12];
assign v__4294_out0 = v_CIN_1159_out0[13:13];
assign v__4327_out0 = v_CIN_1159_out0[14:14];
assign v__5288_out0 = v_CIN_1159_out0[5:5];
assign v__6636_out0 = v_CIN_1159_out0[4:4];
assign v_RM_1809_out0 = v__3768_out0;
assign v_RM_1810_out0 = v__4327_out0;
assign v_RM_1812_out0 = v__5288_out0;
assign v_RM_1813_out0 = v__6636_out0;
assign v_RM_1814_out0 = v__4294_out0;
assign v_RM_1815_out0 = v__1500_out0;
assign v_RM_1816_out0 = v__1893_out0;
assign v_RM_1817_out0 = v__1875_out0;
assign v_RM_1818_out0 = v__1062_out0;
assign v_RM_1819_out0 = v__879_out0;
assign v_RM_1820_out0 = v__1542_out0;
assign v_RM_1821_out0 = v__3352_out0;
assign v_RM_1822_out0 = v__241_out0;
assign v_RM_1823_out0 = v__1516_out0;
assign v_CIN_5014_out0 = v__1081_out0;
assign v_RM_5946_out0 = v__1232_out0;
assign v_RD_3248_out0 = v_CIN_5014_out0;
assign v_G1_4174_out0 = ((v_RD_3255_out0 && !v_RM_5946_out0) || (!v_RD_3255_out0) && v_RM_5946_out0);
assign v_RM_5934_out0 = v_RM_1809_out0;
assign v_RM_5936_out0 = v_RM_1810_out0;
assign v_RM_5940_out0 = v_RM_1812_out0;
assign v_RM_5942_out0 = v_RM_1813_out0;
assign v_RM_5944_out0 = v_RM_1814_out0;
assign v_RM_5947_out0 = v_RM_1815_out0;
assign v_RM_5949_out0 = v_RM_1816_out0;
assign v_RM_5951_out0 = v_RM_1817_out0;
assign v_RM_5953_out0 = v_RM_1818_out0;
assign v_RM_5955_out0 = v_RM_1819_out0;
assign v_RM_5957_out0 = v_RM_1820_out0;
assign v_RM_5959_out0 = v_RM_1821_out0;
assign v_RM_5961_out0 = v_RM_1822_out0;
assign v_RM_5963_out0 = v_RM_1823_out0;
assign v_G2_6419_out0 = v_RD_3255_out0 && v_RM_5946_out0;
assign v_CARRY_2756_out0 = v_G2_6419_out0;
assign v_G1_4162_out0 = ((v_RD_3243_out0 && !v_RM_5934_out0) || (!v_RD_3243_out0) && v_RM_5934_out0);
assign v_G1_4164_out0 = ((v_RD_3245_out0 && !v_RM_5936_out0) || (!v_RD_3245_out0) && v_RM_5936_out0);
assign v_G1_4168_out0 = ((v_RD_3249_out0 && !v_RM_5940_out0) || (!v_RD_3249_out0) && v_RM_5940_out0);
assign v_G1_4170_out0 = ((v_RD_3251_out0 && !v_RM_5942_out0) || (!v_RD_3251_out0) && v_RM_5942_out0);
assign v_G1_4172_out0 = ((v_RD_3253_out0 && !v_RM_5944_out0) || (!v_RD_3253_out0) && v_RM_5944_out0);
assign v_G1_4175_out0 = ((v_RD_3256_out0 && !v_RM_5947_out0) || (!v_RD_3256_out0) && v_RM_5947_out0);
assign v_G1_4177_out0 = ((v_RD_3258_out0 && !v_RM_5949_out0) || (!v_RD_3258_out0) && v_RM_5949_out0);
assign v_G1_4179_out0 = ((v_RD_3260_out0 && !v_RM_5951_out0) || (!v_RD_3260_out0) && v_RM_5951_out0);
assign v_G1_4181_out0 = ((v_RD_3262_out0 && !v_RM_5953_out0) || (!v_RD_3262_out0) && v_RM_5953_out0);
assign v_G1_4183_out0 = ((v_RD_3264_out0 && !v_RM_5955_out0) || (!v_RD_3264_out0) && v_RM_5955_out0);
assign v_G1_4185_out0 = ((v_RD_3266_out0 && !v_RM_5957_out0) || (!v_RD_3266_out0) && v_RM_5957_out0);
assign v_G1_4187_out0 = ((v_RD_3268_out0 && !v_RM_5959_out0) || (!v_RD_3268_out0) && v_RM_5959_out0);
assign v_G1_4189_out0 = ((v_RD_3270_out0 && !v_RM_5961_out0) || (!v_RD_3270_out0) && v_RM_5961_out0);
assign v_G1_4191_out0 = ((v_RD_3272_out0 && !v_RM_5963_out0) || (!v_RD_3272_out0) && v_RM_5963_out0);
assign v_S_4743_out0 = v_G1_4174_out0;
assign v_G2_6407_out0 = v_RD_3243_out0 && v_RM_5934_out0;
assign v_G2_6409_out0 = v_RD_3245_out0 && v_RM_5936_out0;
assign v_G2_6413_out0 = v_RD_3249_out0 && v_RM_5940_out0;
assign v_G2_6415_out0 = v_RD_3251_out0 && v_RM_5942_out0;
assign v_G2_6417_out0 = v_RD_3253_out0 && v_RM_5944_out0;
assign v_G2_6420_out0 = v_RD_3256_out0 && v_RM_5947_out0;
assign v_G2_6422_out0 = v_RD_3258_out0 && v_RM_5949_out0;
assign v_G2_6424_out0 = v_RD_3260_out0 && v_RM_5951_out0;
assign v_G2_6426_out0 = v_RD_3262_out0 && v_RM_5953_out0;
assign v_G2_6428_out0 = v_RD_3264_out0 && v_RM_5955_out0;
assign v_G2_6430_out0 = v_RD_3266_out0 && v_RM_5957_out0;
assign v_G2_6432_out0 = v_RD_3268_out0 && v_RM_5959_out0;
assign v_G2_6434_out0 = v_RD_3270_out0 && v_RM_5961_out0;
assign v_G2_6436_out0 = v_RD_3272_out0 && v_RM_5963_out0;
assign v_S_2290_out0 = v_S_4743_out0;
assign v_CARRY_2744_out0 = v_G2_6407_out0;
assign v_CARRY_2746_out0 = v_G2_6409_out0;
assign v_CARRY_2750_out0 = v_G2_6413_out0;
assign v_CARRY_2752_out0 = v_G2_6415_out0;
assign v_CARRY_2754_out0 = v_G2_6417_out0;
assign v_CARRY_2757_out0 = v_G2_6420_out0;
assign v_CARRY_2759_out0 = v_G2_6422_out0;
assign v_CARRY_2761_out0 = v_G2_6424_out0;
assign v_CARRY_2763_out0 = v_G2_6426_out0;
assign v_CARRY_2765_out0 = v_G2_6428_out0;
assign v_CARRY_2767_out0 = v_G2_6430_out0;
assign v_CARRY_2769_out0 = v_G2_6432_out0;
assign v_CARRY_2771_out0 = v_G2_6434_out0;
assign v_CARRY_2773_out0 = v_G2_6436_out0;
assign v_S_4731_out0 = v_G1_4162_out0;
assign v_S_4733_out0 = v_G1_4164_out0;
assign v_S_4737_out0 = v_G1_4168_out0;
assign v_S_4739_out0 = v_G1_4170_out0;
assign v_S_4741_out0 = v_G1_4172_out0;
assign v_S_4744_out0 = v_G1_4175_out0;
assign v_S_4746_out0 = v_G1_4177_out0;
assign v_S_4748_out0 = v_G1_4179_out0;
assign v_S_4750_out0 = v_G1_4181_out0;
assign v_S_4752_out0 = v_G1_4183_out0;
assign v_S_4754_out0 = v_G1_4185_out0;
assign v_S_4756_out0 = v_G1_4187_out0;
assign v_S_4758_out0 = v_G1_4189_out0;
assign v_S_4760_out0 = v_G1_4191_out0;
assign v_CIN_5020_out0 = v_CARRY_2756_out0;
assign v_RD_3261_out0 = v_CIN_5020_out0;
assign v__5300_out0 = { v__4830_out0,v_S_2290_out0 };
assign v_RM_5935_out0 = v_S_4731_out0;
assign v_RM_5937_out0 = v_S_4733_out0;
assign v_RM_5941_out0 = v_S_4737_out0;
assign v_RM_5943_out0 = v_S_4739_out0;
assign v_RM_5945_out0 = v_S_4741_out0;
assign v_RM_5948_out0 = v_S_4744_out0;
assign v_RM_5950_out0 = v_S_4746_out0;
assign v_RM_5952_out0 = v_S_4748_out0;
assign v_RM_5954_out0 = v_S_4750_out0;
assign v_RM_5956_out0 = v_S_4752_out0;
assign v_RM_5958_out0 = v_S_4754_out0;
assign v_RM_5960_out0 = v_S_4756_out0;
assign v_RM_5962_out0 = v_S_4758_out0;
assign v_RM_5964_out0 = v_S_4760_out0;
assign v_G1_4180_out0 = ((v_RD_3261_out0 && !v_RM_5952_out0) || (!v_RD_3261_out0) && v_RM_5952_out0);
assign v_G2_6425_out0 = v_RD_3261_out0 && v_RM_5952_out0;
assign v_CARRY_2762_out0 = v_G2_6425_out0;
assign v_S_4749_out0 = v_G1_4180_out0;
assign v_S_784_out0 = v_S_4749_out0;
assign v_G1_2136_out0 = v_CARRY_2762_out0 || v_CARRY_2761_out0;
assign v_COUT_520_out0 = v_G1_2136_out0;
assign v_CIN_5026_out0 = v_COUT_520_out0;
assign v_RD_3273_out0 = v_CIN_5026_out0;
assign v_G1_4192_out0 = ((v_RD_3273_out0 && !v_RM_5964_out0) || (!v_RD_3273_out0) && v_RM_5964_out0);
assign v_G2_6437_out0 = v_RD_3273_out0 && v_RM_5964_out0;
assign v_CARRY_2774_out0 = v_G2_6437_out0;
assign v_S_4761_out0 = v_G1_4192_out0;
assign v_S_790_out0 = v_S_4761_out0;
assign v_G1_2142_out0 = v_CARRY_2774_out0 || v_CARRY_2773_out0;
assign v_COUT_526_out0 = v_G1_2142_out0;
assign v__2347_out0 = { v_S_784_out0,v_S_790_out0 };
assign v_CIN_5021_out0 = v_COUT_526_out0;
assign v_RD_3263_out0 = v_CIN_5021_out0;
assign v_G1_4182_out0 = ((v_RD_3263_out0 && !v_RM_5954_out0) || (!v_RD_3263_out0) && v_RM_5954_out0);
assign v_G2_6427_out0 = v_RD_3263_out0 && v_RM_5954_out0;
assign v_CARRY_2764_out0 = v_G2_6427_out0;
assign v_S_4751_out0 = v_G1_4182_out0;
assign v_S_785_out0 = v_S_4751_out0;
assign v_G1_2137_out0 = v_CARRY_2764_out0 || v_CARRY_2763_out0;
assign v_COUT_521_out0 = v_G1_2137_out0;
assign v__1256_out0 = { v__2347_out0,v_S_785_out0 };
assign v_CIN_5016_out0 = v_COUT_521_out0;
assign v_RD_3252_out0 = v_CIN_5016_out0;
assign v_G1_4171_out0 = ((v_RD_3252_out0 && !v_RM_5943_out0) || (!v_RD_3252_out0) && v_RM_5943_out0);
assign v_G2_6416_out0 = v_RD_3252_out0 && v_RM_5943_out0;
assign v_CARRY_2753_out0 = v_G2_6416_out0;
assign v_S_4740_out0 = v_G1_4171_out0;
assign v_S_780_out0 = v_S_4740_out0;
assign v_G1_2132_out0 = v_CARRY_2753_out0 || v_CARRY_2752_out0;
assign v_COUT_516_out0 = v_G1_2132_out0;
assign v__3464_out0 = { v__1256_out0,v_S_780_out0 };
assign v_CIN_5015_out0 = v_COUT_516_out0;
assign v_RD_3250_out0 = v_CIN_5015_out0;
assign v_G1_4169_out0 = ((v_RD_3250_out0 && !v_RM_5941_out0) || (!v_RD_3250_out0) && v_RM_5941_out0);
assign v_G2_6414_out0 = v_RD_3250_out0 && v_RM_5941_out0;
assign v_CARRY_2751_out0 = v_G2_6414_out0;
assign v_S_4738_out0 = v_G1_4169_out0;
assign v_S_779_out0 = v_S_4738_out0;
assign v_G1_2131_out0 = v_CARRY_2751_out0 || v_CARRY_2750_out0;
assign v_COUT_515_out0 = v_G1_2131_out0;
assign v__6674_out0 = { v__3464_out0,v_S_779_out0 };
assign v_CIN_5022_out0 = v_COUT_515_out0;
assign v_RD_3265_out0 = v_CIN_5022_out0;
assign v_G1_4184_out0 = ((v_RD_3265_out0 && !v_RM_5956_out0) || (!v_RD_3265_out0) && v_RM_5956_out0);
assign v_G2_6429_out0 = v_RD_3265_out0 && v_RM_5956_out0;
assign v_CARRY_2766_out0 = v_G2_6429_out0;
assign v_S_4753_out0 = v_G1_4184_out0;
assign v_S_786_out0 = v_S_4753_out0;
assign v_G1_2138_out0 = v_CARRY_2766_out0 || v_CARRY_2765_out0;
assign v_COUT_522_out0 = v_G1_2138_out0;
assign v__1622_out0 = { v__6674_out0,v_S_786_out0 };
assign v_CIN_5023_out0 = v_COUT_522_out0;
assign v_RD_3267_out0 = v_CIN_5023_out0;
assign v_G1_4186_out0 = ((v_RD_3267_out0 && !v_RM_5958_out0) || (!v_RD_3267_out0) && v_RM_5958_out0);
assign v_G2_6431_out0 = v_RD_3267_out0 && v_RM_5958_out0;
assign v_CARRY_2768_out0 = v_G2_6431_out0;
assign v_S_4755_out0 = v_G1_4186_out0;
assign v_S_787_out0 = v_S_4755_out0;
assign v_G1_2139_out0 = v_CARRY_2768_out0 || v_CARRY_2767_out0;
assign v_COUT_523_out0 = v_G1_2139_out0;
assign v__3519_out0 = { v__1622_out0,v_S_787_out0 };
assign v_CIN_5025_out0 = v_COUT_523_out0;
assign v_RD_3271_out0 = v_CIN_5025_out0;
assign v_G1_4190_out0 = ((v_RD_3271_out0 && !v_RM_5962_out0) || (!v_RD_3271_out0) && v_RM_5962_out0);
assign v_G2_6435_out0 = v_RD_3271_out0 && v_RM_5962_out0;
assign v_CARRY_2772_out0 = v_G2_6435_out0;
assign v_S_4759_out0 = v_G1_4190_out0;
assign v_S_789_out0 = v_S_4759_out0;
assign v_G1_2141_out0 = v_CARRY_2772_out0 || v_CARRY_2771_out0;
assign v_COUT_525_out0 = v_G1_2141_out0;
assign v__2330_out0 = { v__3519_out0,v_S_789_out0 };
assign v_CIN_5018_out0 = v_COUT_525_out0;
assign v_RD_3257_out0 = v_CIN_5018_out0;
assign v_G1_4176_out0 = ((v_RD_3257_out0 && !v_RM_5948_out0) || (!v_RD_3257_out0) && v_RM_5948_out0);
assign v_G2_6421_out0 = v_RD_3257_out0 && v_RM_5948_out0;
assign v_CARRY_2758_out0 = v_G2_6421_out0;
assign v_S_4745_out0 = v_G1_4176_out0;
assign v_S_782_out0 = v_S_4745_out0;
assign v_G1_2134_out0 = v_CARRY_2758_out0 || v_CARRY_2757_out0;
assign v_COUT_518_out0 = v_G1_2134_out0;
assign v__3412_out0 = { v__2330_out0,v_S_782_out0 };
assign v_CIN_5019_out0 = v_COUT_518_out0;
assign v_RD_3259_out0 = v_CIN_5019_out0;
assign v_G1_4178_out0 = ((v_RD_3259_out0 && !v_RM_5950_out0) || (!v_RD_3259_out0) && v_RM_5950_out0);
assign v_G2_6423_out0 = v_RD_3259_out0 && v_RM_5950_out0;
assign v_CARRY_2760_out0 = v_G2_6423_out0;
assign v_S_4747_out0 = v_G1_4178_out0;
assign v_S_783_out0 = v_S_4747_out0;
assign v_G1_2135_out0 = v_CARRY_2760_out0 || v_CARRY_2759_out0;
assign v_COUT_519_out0 = v_G1_2135_out0;
assign v__2856_out0 = { v__3412_out0,v_S_783_out0 };
assign v_CIN_5024_out0 = v_COUT_519_out0;
assign v_RD_3269_out0 = v_CIN_5024_out0;
assign v_G1_4188_out0 = ((v_RD_3269_out0 && !v_RM_5960_out0) || (!v_RD_3269_out0) && v_RM_5960_out0);
assign v_G2_6433_out0 = v_RD_3269_out0 && v_RM_5960_out0;
assign v_CARRY_2770_out0 = v_G2_6433_out0;
assign v_S_4757_out0 = v_G1_4188_out0;
assign v_S_788_out0 = v_S_4757_out0;
assign v_G1_2140_out0 = v_CARRY_2770_out0 || v_CARRY_2769_out0;
assign v_COUT_524_out0 = v_G1_2140_out0;
assign v__1000_out0 = { v__2856_out0,v_S_788_out0 };
assign v_CIN_5012_out0 = v_COUT_524_out0;
assign v_RD_3244_out0 = v_CIN_5012_out0;
assign v_G1_4163_out0 = ((v_RD_3244_out0 && !v_RM_5935_out0) || (!v_RD_3244_out0) && v_RM_5935_out0);
assign v_G2_6408_out0 = v_RD_3244_out0 && v_RM_5935_out0;
assign v_CARRY_2745_out0 = v_G2_6408_out0;
assign v_S_4732_out0 = v_G1_4163_out0;
assign v_S_776_out0 = v_S_4732_out0;
assign v_G1_2128_out0 = v_CARRY_2745_out0 || v_CARRY_2744_out0;
assign v_COUT_512_out0 = v_G1_2128_out0;
assign v__1376_out0 = { v__1000_out0,v_S_776_out0 };
assign v_CIN_5017_out0 = v_COUT_512_out0;
assign v_RD_3254_out0 = v_CIN_5017_out0;
assign v_G1_4173_out0 = ((v_RD_3254_out0 && !v_RM_5945_out0) || (!v_RD_3254_out0) && v_RM_5945_out0);
assign v_G2_6418_out0 = v_RD_3254_out0 && v_RM_5945_out0;
assign v_CARRY_2755_out0 = v_G2_6418_out0;
assign v_S_4742_out0 = v_G1_4173_out0;
assign v_S_781_out0 = v_S_4742_out0;
assign v_G1_2133_out0 = v_CARRY_2755_out0 || v_CARRY_2754_out0;
assign v_COUT_517_out0 = v_G1_2133_out0;
assign v__903_out0 = { v__1376_out0,v_S_781_out0 };
assign v_CIN_5013_out0 = v_COUT_517_out0;
assign v_RD_3246_out0 = v_CIN_5013_out0;
assign v_G1_4165_out0 = ((v_RD_3246_out0 && !v_RM_5937_out0) || (!v_RD_3246_out0) && v_RM_5937_out0);
assign v_G2_6410_out0 = v_RD_3246_out0 && v_RM_5937_out0;
assign v_CARRY_2747_out0 = v_G2_6410_out0;
assign v_S_4734_out0 = v_G1_4165_out0;
assign v_S_777_out0 = v_S_4734_out0;
assign v_G1_2129_out0 = v_CARRY_2747_out0 || v_CARRY_2746_out0;
assign v_COUT_513_out0 = v_G1_2129_out0;
assign v__2232_out0 = { v__903_out0,v_S_777_out0 };
assign v_RM_1811_out0 = v_COUT_513_out0;
assign v_RM_5938_out0 = v_RM_1811_out0;
assign v_G1_4166_out0 = ((v_RD_3247_out0 && !v_RM_5938_out0) || (!v_RD_3247_out0) && v_RM_5938_out0);
assign v_G2_6411_out0 = v_RD_3247_out0 && v_RM_5938_out0;
assign v_CARRY_2748_out0 = v_G2_6411_out0;
assign v_S_4735_out0 = v_G1_4166_out0;
assign v_RM_5939_out0 = v_S_4735_out0;
assign v_G1_4167_out0 = ((v_RD_3248_out0 && !v_RM_5939_out0) || (!v_RD_3248_out0) && v_RM_5939_out0);
assign v_G2_6412_out0 = v_RD_3248_out0 && v_RM_5939_out0;
assign v_CARRY_2749_out0 = v_G2_6412_out0;
assign v_S_4736_out0 = v_G1_4167_out0;
assign v_S_778_out0 = v_S_4736_out0;
assign v_G1_2130_out0 = v_CARRY_2749_out0 || v_CARRY_2748_out0;
assign v_COUT_514_out0 = v_G1_2130_out0;
assign v__5255_out0 = { v__2232_out0,v_S_778_out0 };
assign v__5398_out0 = { v__5255_out0,v_COUT_514_out0 };
assign v_COUT_5383_out0 = v__5398_out0;
assign v_CIN_1154_out0 = v_COUT_5383_out0;
assign v__236_out0 = v_CIN_1154_out0[8:8];
assign v__874_out0 = v_CIN_1154_out0[6:6];
assign v__1057_out0 = v_CIN_1154_out0[3:3];
assign v__1076_out0 = v_CIN_1154_out0[15:15];
assign v__1227_out0 = v_CIN_1154_out0[0:0];
assign v__1495_out0 = v_CIN_1154_out0[9:9];
assign v__1511_out0 = v_CIN_1154_out0[2:2];
assign v__1537_out0 = v_CIN_1154_out0[7:7];
assign v__1870_out0 = v_CIN_1154_out0[1:1];
assign v__1888_out0 = v_CIN_1154_out0[10:10];
assign v__3347_out0 = v_CIN_1154_out0[11:11];
assign v__3763_out0 = v_CIN_1154_out0[12:12];
assign v__4289_out0 = v_CIN_1154_out0[13:13];
assign v__4322_out0 = v_CIN_1154_out0[14:14];
assign v__5283_out0 = v_CIN_1154_out0[5:5];
assign v__6631_out0 = v_CIN_1154_out0[4:4];
assign v_RM_1734_out0 = v__3763_out0;
assign v_RM_1735_out0 = v__4322_out0;
assign v_RM_1737_out0 = v__5283_out0;
assign v_RM_1738_out0 = v__6631_out0;
assign v_RM_1739_out0 = v__4289_out0;
assign v_RM_1740_out0 = v__1495_out0;
assign v_RM_1741_out0 = v__1888_out0;
assign v_RM_1742_out0 = v__1870_out0;
assign v_RM_1743_out0 = v__1057_out0;
assign v_RM_1744_out0 = v__874_out0;
assign v_RM_1745_out0 = v__1537_out0;
assign v_RM_1746_out0 = v__3347_out0;
assign v_RM_1747_out0 = v__236_out0;
assign v_RM_1748_out0 = v__1511_out0;
assign v_CIN_4939_out0 = v__1076_out0;
assign v_RM_5791_out0 = v__1227_out0;
assign v_RD_3093_out0 = v_CIN_4939_out0;
assign v_G1_4019_out0 = ((v_RD_3100_out0 && !v_RM_5791_out0) || (!v_RD_3100_out0) && v_RM_5791_out0);
assign v_RM_5779_out0 = v_RM_1734_out0;
assign v_RM_5781_out0 = v_RM_1735_out0;
assign v_RM_5785_out0 = v_RM_1737_out0;
assign v_RM_5787_out0 = v_RM_1738_out0;
assign v_RM_5789_out0 = v_RM_1739_out0;
assign v_RM_5792_out0 = v_RM_1740_out0;
assign v_RM_5794_out0 = v_RM_1741_out0;
assign v_RM_5796_out0 = v_RM_1742_out0;
assign v_RM_5798_out0 = v_RM_1743_out0;
assign v_RM_5800_out0 = v_RM_1744_out0;
assign v_RM_5802_out0 = v_RM_1745_out0;
assign v_RM_5804_out0 = v_RM_1746_out0;
assign v_RM_5806_out0 = v_RM_1747_out0;
assign v_RM_5808_out0 = v_RM_1748_out0;
assign v_G2_6264_out0 = v_RD_3100_out0 && v_RM_5791_out0;
assign v_CARRY_2601_out0 = v_G2_6264_out0;
assign v_G1_4007_out0 = ((v_RD_3088_out0 && !v_RM_5779_out0) || (!v_RD_3088_out0) && v_RM_5779_out0);
assign v_G1_4009_out0 = ((v_RD_3090_out0 && !v_RM_5781_out0) || (!v_RD_3090_out0) && v_RM_5781_out0);
assign v_G1_4013_out0 = ((v_RD_3094_out0 && !v_RM_5785_out0) || (!v_RD_3094_out0) && v_RM_5785_out0);
assign v_G1_4015_out0 = ((v_RD_3096_out0 && !v_RM_5787_out0) || (!v_RD_3096_out0) && v_RM_5787_out0);
assign v_G1_4017_out0 = ((v_RD_3098_out0 && !v_RM_5789_out0) || (!v_RD_3098_out0) && v_RM_5789_out0);
assign v_G1_4020_out0 = ((v_RD_3101_out0 && !v_RM_5792_out0) || (!v_RD_3101_out0) && v_RM_5792_out0);
assign v_G1_4022_out0 = ((v_RD_3103_out0 && !v_RM_5794_out0) || (!v_RD_3103_out0) && v_RM_5794_out0);
assign v_G1_4024_out0 = ((v_RD_3105_out0 && !v_RM_5796_out0) || (!v_RD_3105_out0) && v_RM_5796_out0);
assign v_G1_4026_out0 = ((v_RD_3107_out0 && !v_RM_5798_out0) || (!v_RD_3107_out0) && v_RM_5798_out0);
assign v_G1_4028_out0 = ((v_RD_3109_out0 && !v_RM_5800_out0) || (!v_RD_3109_out0) && v_RM_5800_out0);
assign v_G1_4030_out0 = ((v_RD_3111_out0 && !v_RM_5802_out0) || (!v_RD_3111_out0) && v_RM_5802_out0);
assign v_G1_4032_out0 = ((v_RD_3113_out0 && !v_RM_5804_out0) || (!v_RD_3113_out0) && v_RM_5804_out0);
assign v_G1_4034_out0 = ((v_RD_3115_out0 && !v_RM_5806_out0) || (!v_RD_3115_out0) && v_RM_5806_out0);
assign v_G1_4036_out0 = ((v_RD_3117_out0 && !v_RM_5808_out0) || (!v_RD_3117_out0) && v_RM_5808_out0);
assign v_S_4588_out0 = v_G1_4019_out0;
assign v_G2_6252_out0 = v_RD_3088_out0 && v_RM_5779_out0;
assign v_G2_6254_out0 = v_RD_3090_out0 && v_RM_5781_out0;
assign v_G2_6258_out0 = v_RD_3094_out0 && v_RM_5785_out0;
assign v_G2_6260_out0 = v_RD_3096_out0 && v_RM_5787_out0;
assign v_G2_6262_out0 = v_RD_3098_out0 && v_RM_5789_out0;
assign v_G2_6265_out0 = v_RD_3101_out0 && v_RM_5792_out0;
assign v_G2_6267_out0 = v_RD_3103_out0 && v_RM_5794_out0;
assign v_G2_6269_out0 = v_RD_3105_out0 && v_RM_5796_out0;
assign v_G2_6271_out0 = v_RD_3107_out0 && v_RM_5798_out0;
assign v_G2_6273_out0 = v_RD_3109_out0 && v_RM_5800_out0;
assign v_G2_6275_out0 = v_RD_3111_out0 && v_RM_5802_out0;
assign v_G2_6277_out0 = v_RD_3113_out0 && v_RM_5804_out0;
assign v_G2_6279_out0 = v_RD_3115_out0 && v_RM_5806_out0;
assign v_G2_6281_out0 = v_RD_3117_out0 && v_RM_5808_out0;
assign v_S_2285_out0 = v_S_4588_out0;
assign v_CARRY_2589_out0 = v_G2_6252_out0;
assign v_CARRY_2591_out0 = v_G2_6254_out0;
assign v_CARRY_2595_out0 = v_G2_6258_out0;
assign v_CARRY_2597_out0 = v_G2_6260_out0;
assign v_CARRY_2599_out0 = v_G2_6262_out0;
assign v_CARRY_2602_out0 = v_G2_6265_out0;
assign v_CARRY_2604_out0 = v_G2_6267_out0;
assign v_CARRY_2606_out0 = v_G2_6269_out0;
assign v_CARRY_2608_out0 = v_G2_6271_out0;
assign v_CARRY_2610_out0 = v_G2_6273_out0;
assign v_CARRY_2612_out0 = v_G2_6275_out0;
assign v_CARRY_2614_out0 = v_G2_6277_out0;
assign v_CARRY_2616_out0 = v_G2_6279_out0;
assign v_CARRY_2618_out0 = v_G2_6281_out0;
assign v_S_4576_out0 = v_G1_4007_out0;
assign v_S_4578_out0 = v_G1_4009_out0;
assign v_S_4582_out0 = v_G1_4013_out0;
assign v_S_4584_out0 = v_G1_4015_out0;
assign v_S_4586_out0 = v_G1_4017_out0;
assign v_S_4589_out0 = v_G1_4020_out0;
assign v_S_4591_out0 = v_G1_4022_out0;
assign v_S_4593_out0 = v_G1_4024_out0;
assign v_S_4595_out0 = v_G1_4026_out0;
assign v_S_4597_out0 = v_G1_4028_out0;
assign v_S_4599_out0 = v_G1_4030_out0;
assign v_S_4601_out0 = v_G1_4032_out0;
assign v_S_4603_out0 = v_G1_4034_out0;
assign v_S_4605_out0 = v_G1_4036_out0;
assign v_CIN_4945_out0 = v_CARRY_2601_out0;
assign v_RD_3106_out0 = v_CIN_4945_out0;
assign v_RM_5780_out0 = v_S_4576_out0;
assign v_RM_5782_out0 = v_S_4578_out0;
assign v_RM_5786_out0 = v_S_4582_out0;
assign v_RM_5788_out0 = v_S_4584_out0;
assign v_RM_5790_out0 = v_S_4586_out0;
assign v_RM_5793_out0 = v_S_4589_out0;
assign v_RM_5795_out0 = v_S_4591_out0;
assign v_RM_5797_out0 = v_S_4593_out0;
assign v_RM_5799_out0 = v_S_4595_out0;
assign v_RM_5801_out0 = v_S_4597_out0;
assign v_RM_5803_out0 = v_S_4599_out0;
assign v_RM_5805_out0 = v_S_4601_out0;
assign v_RM_5807_out0 = v_S_4603_out0;
assign v_RM_5809_out0 = v_S_4605_out0;
assign v__6753_out0 = { v__5300_out0,v_S_2285_out0 };
assign v_G1_4025_out0 = ((v_RD_3106_out0 && !v_RM_5797_out0) || (!v_RD_3106_out0) && v_RM_5797_out0);
assign v_G2_6270_out0 = v_RD_3106_out0 && v_RM_5797_out0;
assign v_CARRY_2607_out0 = v_G2_6270_out0;
assign v_S_4594_out0 = v_G1_4025_out0;
assign v_S_709_out0 = v_S_4594_out0;
assign v_G1_2061_out0 = v_CARRY_2607_out0 || v_CARRY_2606_out0;
assign v_COUT_445_out0 = v_G1_2061_out0;
assign v_CIN_4951_out0 = v_COUT_445_out0;
assign v_RD_3118_out0 = v_CIN_4951_out0;
assign v_G1_4037_out0 = ((v_RD_3118_out0 && !v_RM_5809_out0) || (!v_RD_3118_out0) && v_RM_5809_out0);
assign v_G2_6282_out0 = v_RD_3118_out0 && v_RM_5809_out0;
assign v_CARRY_2619_out0 = v_G2_6282_out0;
assign v_S_4606_out0 = v_G1_4037_out0;
assign v_S_715_out0 = v_S_4606_out0;
assign v_G1_2067_out0 = v_CARRY_2619_out0 || v_CARRY_2618_out0;
assign v_COUT_451_out0 = v_G1_2067_out0;
assign v__2342_out0 = { v_S_709_out0,v_S_715_out0 };
assign v_CIN_4946_out0 = v_COUT_451_out0;
assign v_RD_3108_out0 = v_CIN_4946_out0;
assign v_G1_4027_out0 = ((v_RD_3108_out0 && !v_RM_5799_out0) || (!v_RD_3108_out0) && v_RM_5799_out0);
assign v_G2_6272_out0 = v_RD_3108_out0 && v_RM_5799_out0;
assign v_CARRY_2609_out0 = v_G2_6272_out0;
assign v_S_4596_out0 = v_G1_4027_out0;
assign v_S_710_out0 = v_S_4596_out0;
assign v_G1_2062_out0 = v_CARRY_2609_out0 || v_CARRY_2608_out0;
assign v_COUT_446_out0 = v_G1_2062_out0;
assign v__1251_out0 = { v__2342_out0,v_S_710_out0 };
assign v_CIN_4941_out0 = v_COUT_446_out0;
assign v_RD_3097_out0 = v_CIN_4941_out0;
assign v_G1_4016_out0 = ((v_RD_3097_out0 && !v_RM_5788_out0) || (!v_RD_3097_out0) && v_RM_5788_out0);
assign v_G2_6261_out0 = v_RD_3097_out0 && v_RM_5788_out0;
assign v_CARRY_2598_out0 = v_G2_6261_out0;
assign v_S_4585_out0 = v_G1_4016_out0;
assign v_S_705_out0 = v_S_4585_out0;
assign v_G1_2057_out0 = v_CARRY_2598_out0 || v_CARRY_2597_out0;
assign v_COUT_441_out0 = v_G1_2057_out0;
assign v__3459_out0 = { v__1251_out0,v_S_705_out0 };
assign v_CIN_4940_out0 = v_COUT_441_out0;
assign v_RD_3095_out0 = v_CIN_4940_out0;
assign v_G1_4014_out0 = ((v_RD_3095_out0 && !v_RM_5786_out0) || (!v_RD_3095_out0) && v_RM_5786_out0);
assign v_G2_6259_out0 = v_RD_3095_out0 && v_RM_5786_out0;
assign v_CARRY_2596_out0 = v_G2_6259_out0;
assign v_S_4583_out0 = v_G1_4014_out0;
assign v_S_704_out0 = v_S_4583_out0;
assign v_G1_2056_out0 = v_CARRY_2596_out0 || v_CARRY_2595_out0;
assign v_COUT_440_out0 = v_G1_2056_out0;
assign v__6669_out0 = { v__3459_out0,v_S_704_out0 };
assign v_CIN_4947_out0 = v_COUT_440_out0;
assign v_RD_3110_out0 = v_CIN_4947_out0;
assign v_G1_4029_out0 = ((v_RD_3110_out0 && !v_RM_5801_out0) || (!v_RD_3110_out0) && v_RM_5801_out0);
assign v_G2_6274_out0 = v_RD_3110_out0 && v_RM_5801_out0;
assign v_CARRY_2611_out0 = v_G2_6274_out0;
assign v_S_4598_out0 = v_G1_4029_out0;
assign v_S_711_out0 = v_S_4598_out0;
assign v_G1_2063_out0 = v_CARRY_2611_out0 || v_CARRY_2610_out0;
assign v_COUT_447_out0 = v_G1_2063_out0;
assign v__1617_out0 = { v__6669_out0,v_S_711_out0 };
assign v_CIN_4948_out0 = v_COUT_447_out0;
assign v_RD_3112_out0 = v_CIN_4948_out0;
assign v_G1_4031_out0 = ((v_RD_3112_out0 && !v_RM_5803_out0) || (!v_RD_3112_out0) && v_RM_5803_out0);
assign v_G2_6276_out0 = v_RD_3112_out0 && v_RM_5803_out0;
assign v_CARRY_2613_out0 = v_G2_6276_out0;
assign v_S_4600_out0 = v_G1_4031_out0;
assign v_S_712_out0 = v_S_4600_out0;
assign v_G1_2064_out0 = v_CARRY_2613_out0 || v_CARRY_2612_out0;
assign v_COUT_448_out0 = v_G1_2064_out0;
assign v__3514_out0 = { v__1617_out0,v_S_712_out0 };
assign v_CIN_4950_out0 = v_COUT_448_out0;
assign v_RD_3116_out0 = v_CIN_4950_out0;
assign v_G1_4035_out0 = ((v_RD_3116_out0 && !v_RM_5807_out0) || (!v_RD_3116_out0) && v_RM_5807_out0);
assign v_G2_6280_out0 = v_RD_3116_out0 && v_RM_5807_out0;
assign v_CARRY_2617_out0 = v_G2_6280_out0;
assign v_S_4604_out0 = v_G1_4035_out0;
assign v_S_714_out0 = v_S_4604_out0;
assign v_G1_2066_out0 = v_CARRY_2617_out0 || v_CARRY_2616_out0;
assign v_COUT_450_out0 = v_G1_2066_out0;
assign v__2325_out0 = { v__3514_out0,v_S_714_out0 };
assign v_CIN_4943_out0 = v_COUT_450_out0;
assign v_RD_3102_out0 = v_CIN_4943_out0;
assign v_G1_4021_out0 = ((v_RD_3102_out0 && !v_RM_5793_out0) || (!v_RD_3102_out0) && v_RM_5793_out0);
assign v_G2_6266_out0 = v_RD_3102_out0 && v_RM_5793_out0;
assign v_CARRY_2603_out0 = v_G2_6266_out0;
assign v_S_4590_out0 = v_G1_4021_out0;
assign v_S_707_out0 = v_S_4590_out0;
assign v_G1_2059_out0 = v_CARRY_2603_out0 || v_CARRY_2602_out0;
assign v_COUT_443_out0 = v_G1_2059_out0;
assign v__3407_out0 = { v__2325_out0,v_S_707_out0 };
assign v_CIN_4944_out0 = v_COUT_443_out0;
assign v_RD_3104_out0 = v_CIN_4944_out0;
assign v_G1_4023_out0 = ((v_RD_3104_out0 && !v_RM_5795_out0) || (!v_RD_3104_out0) && v_RM_5795_out0);
assign v_G2_6268_out0 = v_RD_3104_out0 && v_RM_5795_out0;
assign v_CARRY_2605_out0 = v_G2_6268_out0;
assign v_S_4592_out0 = v_G1_4023_out0;
assign v_S_708_out0 = v_S_4592_out0;
assign v_G1_2060_out0 = v_CARRY_2605_out0 || v_CARRY_2604_out0;
assign v_COUT_444_out0 = v_G1_2060_out0;
assign v__2851_out0 = { v__3407_out0,v_S_708_out0 };
assign v_CIN_4949_out0 = v_COUT_444_out0;
assign v_RD_3114_out0 = v_CIN_4949_out0;
assign v_G1_4033_out0 = ((v_RD_3114_out0 && !v_RM_5805_out0) || (!v_RD_3114_out0) && v_RM_5805_out0);
assign v_G2_6278_out0 = v_RD_3114_out0 && v_RM_5805_out0;
assign v_CARRY_2615_out0 = v_G2_6278_out0;
assign v_S_4602_out0 = v_G1_4033_out0;
assign v_S_713_out0 = v_S_4602_out0;
assign v_G1_2065_out0 = v_CARRY_2615_out0 || v_CARRY_2614_out0;
assign v_COUT_449_out0 = v_G1_2065_out0;
assign v__995_out0 = { v__2851_out0,v_S_713_out0 };
assign v_CIN_4937_out0 = v_COUT_449_out0;
assign v_RD_3089_out0 = v_CIN_4937_out0;
assign v_G1_4008_out0 = ((v_RD_3089_out0 && !v_RM_5780_out0) || (!v_RD_3089_out0) && v_RM_5780_out0);
assign v_G2_6253_out0 = v_RD_3089_out0 && v_RM_5780_out0;
assign v_CARRY_2590_out0 = v_G2_6253_out0;
assign v_S_4577_out0 = v_G1_4008_out0;
assign v_S_701_out0 = v_S_4577_out0;
assign v_G1_2053_out0 = v_CARRY_2590_out0 || v_CARRY_2589_out0;
assign v_COUT_437_out0 = v_G1_2053_out0;
assign v__1371_out0 = { v__995_out0,v_S_701_out0 };
assign v_CIN_4942_out0 = v_COUT_437_out0;
assign v_RD_3099_out0 = v_CIN_4942_out0;
assign v_G1_4018_out0 = ((v_RD_3099_out0 && !v_RM_5790_out0) || (!v_RD_3099_out0) && v_RM_5790_out0);
assign v_G2_6263_out0 = v_RD_3099_out0 && v_RM_5790_out0;
assign v_CARRY_2600_out0 = v_G2_6263_out0;
assign v_S_4587_out0 = v_G1_4018_out0;
assign v_S_706_out0 = v_S_4587_out0;
assign v_G1_2058_out0 = v_CARRY_2600_out0 || v_CARRY_2599_out0;
assign v_COUT_442_out0 = v_G1_2058_out0;
assign v__898_out0 = { v__1371_out0,v_S_706_out0 };
assign v_CIN_4938_out0 = v_COUT_442_out0;
assign v_RD_3091_out0 = v_CIN_4938_out0;
assign v_G1_4010_out0 = ((v_RD_3091_out0 && !v_RM_5782_out0) || (!v_RD_3091_out0) && v_RM_5782_out0);
assign v_G2_6255_out0 = v_RD_3091_out0 && v_RM_5782_out0;
assign v_CARRY_2592_out0 = v_G2_6255_out0;
assign v_S_4579_out0 = v_G1_4010_out0;
assign v_S_702_out0 = v_S_4579_out0;
assign v_G1_2054_out0 = v_CARRY_2592_out0 || v_CARRY_2591_out0;
assign v_COUT_438_out0 = v_G1_2054_out0;
assign v__2227_out0 = { v__898_out0,v_S_702_out0 };
assign v_RM_1736_out0 = v_COUT_438_out0;
assign v_RM_5783_out0 = v_RM_1736_out0;
assign v_G1_4011_out0 = ((v_RD_3092_out0 && !v_RM_5783_out0) || (!v_RD_3092_out0) && v_RM_5783_out0);
assign v_G2_6256_out0 = v_RD_3092_out0 && v_RM_5783_out0;
assign v_CARRY_2593_out0 = v_G2_6256_out0;
assign v_S_4580_out0 = v_G1_4011_out0;
assign v_RM_5784_out0 = v_S_4580_out0;
assign v_G1_4012_out0 = ((v_RD_3093_out0 && !v_RM_5784_out0) || (!v_RD_3093_out0) && v_RM_5784_out0);
assign v_G2_6257_out0 = v_RD_3093_out0 && v_RM_5784_out0;
assign v_CARRY_2594_out0 = v_G2_6257_out0;
assign v_S_4581_out0 = v_G1_4012_out0;
assign v_S_703_out0 = v_S_4581_out0;
assign v_G1_2055_out0 = v_CARRY_2594_out0 || v_CARRY_2593_out0;
assign v_COUT_439_out0 = v_G1_2055_out0;
assign v__5250_out0 = { v__2227_out0,v_S_703_out0 };
assign v__5393_out0 = { v__5250_out0,v_COUT_439_out0 };
assign v_COUT_5378_out0 = v__5393_out0;
assign v_CIN_1153_out0 = v_COUT_5378_out0;
assign v__235_out0 = v_CIN_1153_out0[8:8];
assign v__873_out0 = v_CIN_1153_out0[6:6];
assign v__1056_out0 = v_CIN_1153_out0[3:3];
assign v__1075_out0 = v_CIN_1153_out0[15:15];
assign v__1226_out0 = v_CIN_1153_out0[0:0];
assign v__1494_out0 = v_CIN_1153_out0[9:9];
assign v__1510_out0 = v_CIN_1153_out0[2:2];
assign v__1536_out0 = v_CIN_1153_out0[7:7];
assign v__1869_out0 = v_CIN_1153_out0[1:1];
assign v__1887_out0 = v_CIN_1153_out0[10:10];
assign v__3346_out0 = v_CIN_1153_out0[11:11];
assign v__3762_out0 = v_CIN_1153_out0[12:12];
assign v__4288_out0 = v_CIN_1153_out0[13:13];
assign v__4321_out0 = v_CIN_1153_out0[14:14];
assign v__5282_out0 = v_CIN_1153_out0[5:5];
assign v__6630_out0 = v_CIN_1153_out0[4:4];
assign v_RM_1719_out0 = v__3762_out0;
assign v_RM_1720_out0 = v__4321_out0;
assign v_RM_1722_out0 = v__5282_out0;
assign v_RM_1723_out0 = v__6630_out0;
assign v_RM_1724_out0 = v__4288_out0;
assign v_RM_1725_out0 = v__1494_out0;
assign v_RM_1726_out0 = v__1887_out0;
assign v_RM_1727_out0 = v__1869_out0;
assign v_RM_1728_out0 = v__1056_out0;
assign v_RM_1729_out0 = v__873_out0;
assign v_RM_1730_out0 = v__1536_out0;
assign v_RM_1731_out0 = v__3346_out0;
assign v_RM_1732_out0 = v__235_out0;
assign v_RM_1733_out0 = v__1510_out0;
assign v_CIN_4924_out0 = v__1075_out0;
assign v_RM_5760_out0 = v__1226_out0;
assign v_RD_3062_out0 = v_CIN_4924_out0;
assign v_G1_3988_out0 = ((v_RD_3069_out0 && !v_RM_5760_out0) || (!v_RD_3069_out0) && v_RM_5760_out0);
assign v_RM_5748_out0 = v_RM_1719_out0;
assign v_RM_5750_out0 = v_RM_1720_out0;
assign v_RM_5754_out0 = v_RM_1722_out0;
assign v_RM_5756_out0 = v_RM_1723_out0;
assign v_RM_5758_out0 = v_RM_1724_out0;
assign v_RM_5761_out0 = v_RM_1725_out0;
assign v_RM_5763_out0 = v_RM_1726_out0;
assign v_RM_5765_out0 = v_RM_1727_out0;
assign v_RM_5767_out0 = v_RM_1728_out0;
assign v_RM_5769_out0 = v_RM_1729_out0;
assign v_RM_5771_out0 = v_RM_1730_out0;
assign v_RM_5773_out0 = v_RM_1731_out0;
assign v_RM_5775_out0 = v_RM_1732_out0;
assign v_RM_5777_out0 = v_RM_1733_out0;
assign v_G2_6233_out0 = v_RD_3069_out0 && v_RM_5760_out0;
assign v_CARRY_2570_out0 = v_G2_6233_out0;
assign v_G1_3976_out0 = ((v_RD_3057_out0 && !v_RM_5748_out0) || (!v_RD_3057_out0) && v_RM_5748_out0);
assign v_G1_3978_out0 = ((v_RD_3059_out0 && !v_RM_5750_out0) || (!v_RD_3059_out0) && v_RM_5750_out0);
assign v_G1_3982_out0 = ((v_RD_3063_out0 && !v_RM_5754_out0) || (!v_RD_3063_out0) && v_RM_5754_out0);
assign v_G1_3984_out0 = ((v_RD_3065_out0 && !v_RM_5756_out0) || (!v_RD_3065_out0) && v_RM_5756_out0);
assign v_G1_3986_out0 = ((v_RD_3067_out0 && !v_RM_5758_out0) || (!v_RD_3067_out0) && v_RM_5758_out0);
assign v_G1_3989_out0 = ((v_RD_3070_out0 && !v_RM_5761_out0) || (!v_RD_3070_out0) && v_RM_5761_out0);
assign v_G1_3991_out0 = ((v_RD_3072_out0 && !v_RM_5763_out0) || (!v_RD_3072_out0) && v_RM_5763_out0);
assign v_G1_3993_out0 = ((v_RD_3074_out0 && !v_RM_5765_out0) || (!v_RD_3074_out0) && v_RM_5765_out0);
assign v_G1_3995_out0 = ((v_RD_3076_out0 && !v_RM_5767_out0) || (!v_RD_3076_out0) && v_RM_5767_out0);
assign v_G1_3997_out0 = ((v_RD_3078_out0 && !v_RM_5769_out0) || (!v_RD_3078_out0) && v_RM_5769_out0);
assign v_G1_3999_out0 = ((v_RD_3080_out0 && !v_RM_5771_out0) || (!v_RD_3080_out0) && v_RM_5771_out0);
assign v_G1_4001_out0 = ((v_RD_3082_out0 && !v_RM_5773_out0) || (!v_RD_3082_out0) && v_RM_5773_out0);
assign v_G1_4003_out0 = ((v_RD_3084_out0 && !v_RM_5775_out0) || (!v_RD_3084_out0) && v_RM_5775_out0);
assign v_G1_4005_out0 = ((v_RD_3086_out0 && !v_RM_5777_out0) || (!v_RD_3086_out0) && v_RM_5777_out0);
assign v_S_4557_out0 = v_G1_3988_out0;
assign v_G2_6221_out0 = v_RD_3057_out0 && v_RM_5748_out0;
assign v_G2_6223_out0 = v_RD_3059_out0 && v_RM_5750_out0;
assign v_G2_6227_out0 = v_RD_3063_out0 && v_RM_5754_out0;
assign v_G2_6229_out0 = v_RD_3065_out0 && v_RM_5756_out0;
assign v_G2_6231_out0 = v_RD_3067_out0 && v_RM_5758_out0;
assign v_G2_6234_out0 = v_RD_3070_out0 && v_RM_5761_out0;
assign v_G2_6236_out0 = v_RD_3072_out0 && v_RM_5763_out0;
assign v_G2_6238_out0 = v_RD_3074_out0 && v_RM_5765_out0;
assign v_G2_6240_out0 = v_RD_3076_out0 && v_RM_5767_out0;
assign v_G2_6242_out0 = v_RD_3078_out0 && v_RM_5769_out0;
assign v_G2_6244_out0 = v_RD_3080_out0 && v_RM_5771_out0;
assign v_G2_6246_out0 = v_RD_3082_out0 && v_RM_5773_out0;
assign v_G2_6248_out0 = v_RD_3084_out0 && v_RM_5775_out0;
assign v_G2_6250_out0 = v_RD_3086_out0 && v_RM_5777_out0;
assign v_S_2284_out0 = v_S_4557_out0;
assign v_CARRY_2558_out0 = v_G2_6221_out0;
assign v_CARRY_2560_out0 = v_G2_6223_out0;
assign v_CARRY_2564_out0 = v_G2_6227_out0;
assign v_CARRY_2566_out0 = v_G2_6229_out0;
assign v_CARRY_2568_out0 = v_G2_6231_out0;
assign v_CARRY_2571_out0 = v_G2_6234_out0;
assign v_CARRY_2573_out0 = v_G2_6236_out0;
assign v_CARRY_2575_out0 = v_G2_6238_out0;
assign v_CARRY_2577_out0 = v_G2_6240_out0;
assign v_CARRY_2579_out0 = v_G2_6242_out0;
assign v_CARRY_2581_out0 = v_G2_6244_out0;
assign v_CARRY_2583_out0 = v_G2_6246_out0;
assign v_CARRY_2585_out0 = v_G2_6248_out0;
assign v_CARRY_2587_out0 = v_G2_6250_out0;
assign v_S_4545_out0 = v_G1_3976_out0;
assign v_S_4547_out0 = v_G1_3978_out0;
assign v_S_4551_out0 = v_G1_3982_out0;
assign v_S_4553_out0 = v_G1_3984_out0;
assign v_S_4555_out0 = v_G1_3986_out0;
assign v_S_4558_out0 = v_G1_3989_out0;
assign v_S_4560_out0 = v_G1_3991_out0;
assign v_S_4562_out0 = v_G1_3993_out0;
assign v_S_4564_out0 = v_G1_3995_out0;
assign v_S_4566_out0 = v_G1_3997_out0;
assign v_S_4568_out0 = v_G1_3999_out0;
assign v_S_4570_out0 = v_G1_4001_out0;
assign v_S_4572_out0 = v_G1_4003_out0;
assign v_S_4574_out0 = v_G1_4005_out0;
assign v_CIN_4930_out0 = v_CARRY_2570_out0;
assign v__195_out0 = { v__6753_out0,v_S_2284_out0 };
assign v_RD_3075_out0 = v_CIN_4930_out0;
assign v_RM_5749_out0 = v_S_4545_out0;
assign v_RM_5751_out0 = v_S_4547_out0;
assign v_RM_5755_out0 = v_S_4551_out0;
assign v_RM_5757_out0 = v_S_4553_out0;
assign v_RM_5759_out0 = v_S_4555_out0;
assign v_RM_5762_out0 = v_S_4558_out0;
assign v_RM_5764_out0 = v_S_4560_out0;
assign v_RM_5766_out0 = v_S_4562_out0;
assign v_RM_5768_out0 = v_S_4564_out0;
assign v_RM_5770_out0 = v_S_4566_out0;
assign v_RM_5772_out0 = v_S_4568_out0;
assign v_RM_5774_out0 = v_S_4570_out0;
assign v_RM_5776_out0 = v_S_4572_out0;
assign v_RM_5778_out0 = v_S_4574_out0;
assign v_MUX1_1326_out0 = v_EXEC2_1578_out0 ? v_REG1_6571_out0 : v__195_out0;
assign v_G1_3994_out0 = ((v_RD_3075_out0 && !v_RM_5766_out0) || (!v_RD_3075_out0) && v_RM_5766_out0);
assign v_G2_6239_out0 = v_RD_3075_out0 && v_RM_5766_out0;
assign v_M_REGIN_135_out0 = v_MUX1_1326_out0;
assign v_CARRY_2576_out0 = v_G2_6239_out0;
assign v_S_4563_out0 = v_G1_3994_out0;
assign v_S_694_out0 = v_S_4563_out0;
assign v_MULTI_REGIN_1399_out0 = v_M_REGIN_135_out0;
assign v_G1_2046_out0 = v_CARRY_2576_out0 || v_CARRY_2575_out0;
assign v_COUT_430_out0 = v_G1_2046_out0;
assign v_MULTI_OUT_6706_out0 = v_MULTI_REGIN_1399_out0;
assign v_MULTI_OUT_1589_out0 = v_MULTI_OUT_6706_out0;
assign v_CIN_4936_out0 = v_COUT_430_out0;
assign v_RD_3087_out0 = v_CIN_4936_out0;
assign v_G1_4006_out0 = ((v_RD_3087_out0 && !v_RM_5778_out0) || (!v_RD_3087_out0) && v_RM_5778_out0);
assign v_G2_6251_out0 = v_RD_3087_out0 && v_RM_5778_out0;
assign v_CARRY_2588_out0 = v_G2_6251_out0;
assign v_S_4575_out0 = v_G1_4006_out0;
assign v_S_700_out0 = v_S_4575_out0;
assign v_G1_2052_out0 = v_CARRY_2588_out0 || v_CARRY_2587_out0;
assign v_COUT_436_out0 = v_G1_2052_out0;
assign v__2341_out0 = { v_S_694_out0,v_S_700_out0 };
assign v_CIN_4931_out0 = v_COUT_436_out0;
assign v_RD_3077_out0 = v_CIN_4931_out0;
assign v_G1_3996_out0 = ((v_RD_3077_out0 && !v_RM_5768_out0) || (!v_RD_3077_out0) && v_RM_5768_out0);
assign v_G2_6241_out0 = v_RD_3077_out0 && v_RM_5768_out0;
assign v_CARRY_2578_out0 = v_G2_6241_out0;
assign v_S_4565_out0 = v_G1_3996_out0;
assign v_S_695_out0 = v_S_4565_out0;
assign v_G1_2047_out0 = v_CARRY_2578_out0 || v_CARRY_2577_out0;
assign v_COUT_431_out0 = v_G1_2047_out0;
assign v__1250_out0 = { v__2341_out0,v_S_695_out0 };
assign v_CIN_4926_out0 = v_COUT_431_out0;
assign v_RD_3066_out0 = v_CIN_4926_out0;
assign v_G1_3985_out0 = ((v_RD_3066_out0 && !v_RM_5757_out0) || (!v_RD_3066_out0) && v_RM_5757_out0);
assign v_G2_6230_out0 = v_RD_3066_out0 && v_RM_5757_out0;
assign v_CARRY_2567_out0 = v_G2_6230_out0;
assign v_S_4554_out0 = v_G1_3985_out0;
assign v_S_690_out0 = v_S_4554_out0;
assign v_G1_2042_out0 = v_CARRY_2567_out0 || v_CARRY_2566_out0;
assign v_COUT_426_out0 = v_G1_2042_out0;
assign v__3458_out0 = { v__1250_out0,v_S_690_out0 };
assign v_CIN_4925_out0 = v_COUT_426_out0;
assign v_RD_3064_out0 = v_CIN_4925_out0;
assign v_G1_3983_out0 = ((v_RD_3064_out0 && !v_RM_5755_out0) || (!v_RD_3064_out0) && v_RM_5755_out0);
assign v_G2_6228_out0 = v_RD_3064_out0 && v_RM_5755_out0;
assign v_CARRY_2565_out0 = v_G2_6228_out0;
assign v_S_4552_out0 = v_G1_3983_out0;
assign v_S_689_out0 = v_S_4552_out0;
assign v_G1_2041_out0 = v_CARRY_2565_out0 || v_CARRY_2564_out0;
assign v_COUT_425_out0 = v_G1_2041_out0;
assign v__6668_out0 = { v__3458_out0,v_S_689_out0 };
assign v_CIN_4932_out0 = v_COUT_425_out0;
assign v_RD_3079_out0 = v_CIN_4932_out0;
assign v_G1_3998_out0 = ((v_RD_3079_out0 && !v_RM_5770_out0) || (!v_RD_3079_out0) && v_RM_5770_out0);
assign v_G2_6243_out0 = v_RD_3079_out0 && v_RM_5770_out0;
assign v_CARRY_2580_out0 = v_G2_6243_out0;
assign v_S_4567_out0 = v_G1_3998_out0;
assign v_S_696_out0 = v_S_4567_out0;
assign v_G1_2048_out0 = v_CARRY_2580_out0 || v_CARRY_2579_out0;
assign v_COUT_432_out0 = v_G1_2048_out0;
assign v__1616_out0 = { v__6668_out0,v_S_696_out0 };
assign v_CIN_4933_out0 = v_COUT_432_out0;
assign v_RD_3081_out0 = v_CIN_4933_out0;
assign v_G1_4000_out0 = ((v_RD_3081_out0 && !v_RM_5772_out0) || (!v_RD_3081_out0) && v_RM_5772_out0);
assign v_G2_6245_out0 = v_RD_3081_out0 && v_RM_5772_out0;
assign v_CARRY_2582_out0 = v_G2_6245_out0;
assign v_S_4569_out0 = v_G1_4000_out0;
assign v_S_697_out0 = v_S_4569_out0;
assign v_G1_2049_out0 = v_CARRY_2582_out0 || v_CARRY_2581_out0;
assign v_COUT_433_out0 = v_G1_2049_out0;
assign v__3513_out0 = { v__1616_out0,v_S_697_out0 };
assign v_CIN_4935_out0 = v_COUT_433_out0;
assign v_RD_3085_out0 = v_CIN_4935_out0;
assign v_G1_4004_out0 = ((v_RD_3085_out0 && !v_RM_5776_out0) || (!v_RD_3085_out0) && v_RM_5776_out0);
assign v_G2_6249_out0 = v_RD_3085_out0 && v_RM_5776_out0;
assign v_CARRY_2586_out0 = v_G2_6249_out0;
assign v_S_4573_out0 = v_G1_4004_out0;
assign v_S_699_out0 = v_S_4573_out0;
assign v_G1_2051_out0 = v_CARRY_2586_out0 || v_CARRY_2585_out0;
assign v_COUT_435_out0 = v_G1_2051_out0;
assign v__2324_out0 = { v__3513_out0,v_S_699_out0 };
assign v_CIN_4928_out0 = v_COUT_435_out0;
assign v_RD_3071_out0 = v_CIN_4928_out0;
assign v_G1_3990_out0 = ((v_RD_3071_out0 && !v_RM_5762_out0) || (!v_RD_3071_out0) && v_RM_5762_out0);
assign v_G2_6235_out0 = v_RD_3071_out0 && v_RM_5762_out0;
assign v_CARRY_2572_out0 = v_G2_6235_out0;
assign v_S_4559_out0 = v_G1_3990_out0;
assign v_S_692_out0 = v_S_4559_out0;
assign v_G1_2044_out0 = v_CARRY_2572_out0 || v_CARRY_2571_out0;
assign v_COUT_428_out0 = v_G1_2044_out0;
assign v__3406_out0 = { v__2324_out0,v_S_692_out0 };
assign v_CIN_4929_out0 = v_COUT_428_out0;
assign v_RD_3073_out0 = v_CIN_4929_out0;
assign v_G1_3992_out0 = ((v_RD_3073_out0 && !v_RM_5764_out0) || (!v_RD_3073_out0) && v_RM_5764_out0);
assign v_G2_6237_out0 = v_RD_3073_out0 && v_RM_5764_out0;
assign v_CARRY_2574_out0 = v_G2_6237_out0;
assign v_S_4561_out0 = v_G1_3992_out0;
assign v_S_693_out0 = v_S_4561_out0;
assign v_G1_2045_out0 = v_CARRY_2574_out0 || v_CARRY_2573_out0;
assign v_COUT_429_out0 = v_G1_2045_out0;
assign v__2850_out0 = { v__3406_out0,v_S_693_out0 };
assign v_CIN_4934_out0 = v_COUT_429_out0;
assign v_RD_3083_out0 = v_CIN_4934_out0;
assign v_G1_4002_out0 = ((v_RD_3083_out0 && !v_RM_5774_out0) || (!v_RD_3083_out0) && v_RM_5774_out0);
assign v_G2_6247_out0 = v_RD_3083_out0 && v_RM_5774_out0;
assign v_CARRY_2584_out0 = v_G2_6247_out0;
assign v_S_4571_out0 = v_G1_4002_out0;
assign v_S_698_out0 = v_S_4571_out0;
assign v_G1_2050_out0 = v_CARRY_2584_out0 || v_CARRY_2583_out0;
assign v_COUT_434_out0 = v_G1_2050_out0;
assign v__994_out0 = { v__2850_out0,v_S_698_out0 };
assign v_CIN_4922_out0 = v_COUT_434_out0;
assign v_RD_3058_out0 = v_CIN_4922_out0;
assign v_G1_3977_out0 = ((v_RD_3058_out0 && !v_RM_5749_out0) || (!v_RD_3058_out0) && v_RM_5749_out0);
assign v_G2_6222_out0 = v_RD_3058_out0 && v_RM_5749_out0;
assign v_CARRY_2559_out0 = v_G2_6222_out0;
assign v_S_4546_out0 = v_G1_3977_out0;
assign v_S_686_out0 = v_S_4546_out0;
assign v_G1_2038_out0 = v_CARRY_2559_out0 || v_CARRY_2558_out0;
assign v_COUT_422_out0 = v_G1_2038_out0;
assign v__1370_out0 = { v__994_out0,v_S_686_out0 };
assign v_CIN_4927_out0 = v_COUT_422_out0;
assign v_RD_3068_out0 = v_CIN_4927_out0;
assign v_G1_3987_out0 = ((v_RD_3068_out0 && !v_RM_5759_out0) || (!v_RD_3068_out0) && v_RM_5759_out0);
assign v_G2_6232_out0 = v_RD_3068_out0 && v_RM_5759_out0;
assign v_CARRY_2569_out0 = v_G2_6232_out0;
assign v_S_4556_out0 = v_G1_3987_out0;
assign v_S_691_out0 = v_S_4556_out0;
assign v_G1_2043_out0 = v_CARRY_2569_out0 || v_CARRY_2568_out0;
assign v_COUT_427_out0 = v_G1_2043_out0;
assign v__897_out0 = { v__1370_out0,v_S_691_out0 };
assign v_CIN_4923_out0 = v_COUT_427_out0;
assign v_RD_3060_out0 = v_CIN_4923_out0;
assign v_G1_3979_out0 = ((v_RD_3060_out0 && !v_RM_5751_out0) || (!v_RD_3060_out0) && v_RM_5751_out0);
assign v_G2_6224_out0 = v_RD_3060_out0 && v_RM_5751_out0;
assign v_CARRY_2561_out0 = v_G2_6224_out0;
assign v_S_4548_out0 = v_G1_3979_out0;
assign v_S_687_out0 = v_S_4548_out0;
assign v_G1_2039_out0 = v_CARRY_2561_out0 || v_CARRY_2560_out0;
assign v_COUT_423_out0 = v_G1_2039_out0;
assign v__2226_out0 = { v__897_out0,v_S_687_out0 };
assign v_RM_1721_out0 = v_COUT_423_out0;
assign v_RM_5752_out0 = v_RM_1721_out0;
assign v_G1_3980_out0 = ((v_RD_3061_out0 && !v_RM_5752_out0) || (!v_RD_3061_out0) && v_RM_5752_out0);
assign v_G2_6225_out0 = v_RD_3061_out0 && v_RM_5752_out0;
assign v_CARRY_2562_out0 = v_G2_6225_out0;
assign v_S_4549_out0 = v_G1_3980_out0;
assign v_RM_5753_out0 = v_S_4549_out0;
assign v_G1_3981_out0 = ((v_RD_3062_out0 && !v_RM_5753_out0) || (!v_RD_3062_out0) && v_RM_5753_out0);
assign v_G2_6226_out0 = v_RD_3062_out0 && v_RM_5753_out0;
assign v_CARRY_2563_out0 = v_G2_6226_out0;
assign v_S_4550_out0 = v_G1_3981_out0;
assign v_S_688_out0 = v_S_4550_out0;
assign v_G1_2040_out0 = v_CARRY_2563_out0 || v_CARRY_2562_out0;
assign v_COUT_424_out0 = v_G1_2040_out0;
assign v__5249_out0 = { v__2226_out0,v_S_688_out0 };
assign v__5392_out0 = { v__5249_out0,v_COUT_424_out0 };
assign v_COUT_5377_out0 = v__5392_out0;
assign v__106_out0 = { v__195_out0,v_COUT_5377_out0 };
assign v_FLOATING_MULTI_3782_out0 = v__106_out0;
assign v_32BIT_MULTI_580_out0 = v_FLOATING_MULTI_3782_out0;
assign v_32BITPRODUCT_44_out0 = v_32BIT_MULTI_580_out0;
assign v_32BITPRODUCT_6034_out0 = v_32BITPRODUCT_44_out0;
assign v_SEL7_2367_out0 = v_32BITPRODUCT_6034_out0[21:10];
assign v_MULTI_PRODUCT_3485_out0 = v_SEL7_2367_out0;
assign v_MUX8_6790_out0 = v_MULTI_INSTRUCTION_1193_out0 ? v_MULTI_PRODUCT_3485_out0 : v_SEL8_5260_out0;
assign v_SEL3_561_out0 = v_MUX8_6790_out0[11:11];
assign v_SEL5_1487_out0 = v_MUX8_6790_out0[10:10];
assign v_SEL2_6650_out0 = v_MUX8_6790_out0[10:0];
assign v_SEL6_1948_out0 = v_SEL2_6650_out0[8:0];
assign v_BIT10_3441_out0 = v_SEL5_1487_out0;
assign v_OVERFLOW_5165_out0 = v_SEL3_561_out0;
assign v_SEL4_5525_out0 = v_SEL2_6650_out0[9:0];
assign v_SEL9_6774_out0 = v_SEL2_6650_out0[10:1];
assign v_G3_1313_out0 = v_BIT10_3441_out0 || v_OVERFLOW_5165_out0;
assign v__4272_out0 = { v_C9_1477_out0,v_SEL6_1948_out0 };
assign v_MUX5_5060_out0 = v_SUBNORMAL_4335_out0 ? v_BIT10_3441_out0 : v_OVERFLOW_5165_out0;
assign v_MUX4_5103_out0 = v_OVERFLOW_5165_out0 ? v_SEL9_6774_out0 : v_SEL4_5525_out0;
assign v_G2_2863_out0 = !(v_G3_1313_out0 || v_SUBNORMAL_4335_out0);
assign v_UNDERFLOW_3395_out0 = v_G2_2863_out0;
assign v_G4_1575_out0 = v_UNDERFLOW_3395_out0 && v_G5_309_out0;
assign v_MUX7_2189_out0 = v_UNDERFLOW_3395_out0 ? v_C10_5536_out0 : v_C8_1346_out0;
assign {v_A7_1328_out1,v_A7_1328_out0 } = v_EXP_1188_out0 + v_MUX7_2189_out0 + v_MUX5_5060_out0;
assign v_MUX6_5100_out0 = v_G4_1575_out0 ? v__4272_out0 : v_MUX4_5103_out0;
assign v_SIG_ANS_213_out0 = v_MUX6_5100_out0;
assign v_NOTUSED3_5192_out0 = v_A7_1328_out1;
assign v_EXP_ANS_6772_out0 = v_A7_1328_out0;
assign v_EXP_ANS_981_out0 = v_EXP_ANS_6772_out0;
assign v_SIG_ANS_1139_out0 = v_SIG_ANS_213_out0;
assign v__1272_out0 = { v_EXP_ANS_981_out0,v_SIGN_ANS_4257_out0 };
assign v_SIG_ANS_1593_out0 = v_SIG_ANS_1139_out0;
assign v_EXP_ANS_5163_out0 = v_EXP_ANS_981_out0;
assign v_SIG_ANS_5077_out0 = v_SIG_ANS_1593_out0;
assign v__5146_out0 = { v_SIG_ANS_1139_out0,v__1272_out0 };
assign v_EXP_ANS_5443_out0 = v_EXP_ANS_5163_out0;
assign v_16BIT_WORD_ANSWER_4340_out0 = v__5146_out0;
assign v_FLOATING_REGISTER_IN_275_out0 = v_16BIT_WORD_ANSWER_4340_out0;
assign v_MUX12_840_out0 = v_FLOATING_EN_ALU_307_out0 ? v_FLOATING_REGISTER_IN_275_out0 : v_ALUOUT_2249_out0;
assign v_MUX5_1270_out0 = v_FLOATING_INS_6796_out0 ? v_FLOATING_REGISTER_IN_275_out0 : v_MULTI_REGIN_1399_out0;
assign v_MUX4_6_out0 = v_MULTI_OPCODE_1474_out0 ? v_MUX5_1270_out0 : v_LS_REGIN_1606_out0;
assign v_MUX11_6771_out0 = v_IR15_1201_out0 ? v_MUX12_840_out0 : v_MUX4_6_out0;
assign v_DIN_1105_out0 = v_MUX11_6771_out0;
assign v_DIN3_5083_out0 = v_MUX11_6771_out0;
assign v_DIN_4828_out0 = v_DIN_1105_out0;


endmodule
